// removed module with interface ports: VX_opc_unit
// removed module with interface ports: VX_schedule
module VX_serial_div (
	clk,
	reset,
	strobe,
	busy,
	is_signed,
	numer,
	denom,
	quotient,
	remainder
);
	// Trace: src/VX_serial_div.sv:2:15
	parameter WIDTHN = 32;
	// Trace: src/VX_serial_div.sv:3:15
	parameter WIDTHD = 32;
	// Trace: src/VX_serial_div.sv:4:15
	parameter WIDTHQ = 32;
	// Trace: src/VX_serial_div.sv:5:15
	parameter WIDTHR = 32;
	// Trace: src/VX_serial_div.sv:6:15
	parameter LANES = 1;
	// Trace: src/VX_serial_div.sv:8:5
	input wire clk;
	// Trace: src/VX_serial_div.sv:9:5
	input wire reset;
	// Trace: src/VX_serial_div.sv:10:5
	input wire strobe;
	// Trace: src/VX_serial_div.sv:11:5
	output wire busy;
	// Trace: src/VX_serial_div.sv:12:5
	input wire is_signed;
	// Trace: src/VX_serial_div.sv:13:5
	input wire [(LANES * WIDTHN) - 1:0] numer;
	// Trace: src/VX_serial_div.sv:14:5
	input wire [(LANES * WIDTHD) - 1:0] denom;
	// Trace: src/VX_serial_div.sv:15:5
	output wire [(LANES * WIDTHQ) - 1:0] quotient;
	// Trace: src/VX_serial_div.sv:16:5
	output wire [(LANES * WIDTHR) - 1:0] remainder;
	// Trace: src/VX_serial_div.sv:18:5
	localparam MIN_ND = (WIDTHN < WIDTHD ? WIDTHN : WIDTHD);
	// Trace: src/VX_serial_div.sv:19:5
	localparam CNTRW = $clog2(WIDTHN);
	// Trace: src/VX_serial_div.sv:20:5
	reg [((WIDTHN + MIN_ND) >= 0 ? (LANES * ((WIDTHN + MIN_ND) + 1)) - 1 : (LANES * (1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) - 1)):((WIDTHN + MIN_ND) >= 0 ? 0 : (WIDTHN + MIN_ND) + 0)] working;
	// Trace: src/VX_serial_div.sv:21:5
	reg [(LANES * WIDTHD) - 1:0] denom_r;
	// Trace: src/VX_serial_div.sv:22:5
	wire [(LANES * WIDTHN) - 1:0] numer_qual;
	// Trace: src/VX_serial_div.sv:23:5
	wire [(LANES * WIDTHD) - 1:0] denom_qual;
	// Trace: src/VX_serial_div.sv:24:5
	wire [(WIDTHD >= 0 ? (LANES * (WIDTHD + 1)) - 1 : (LANES * (1 - WIDTHD)) + (WIDTHD - 1)):(WIDTHD >= 0 ? 0 : WIDTHD + 0)] sub_result;
	// Trace: src/VX_serial_div.sv:25:5
	reg [LANES - 1:0] inv_quot;
	reg [LANES - 1:0] inv_rem;
	// Trace: src/VX_serial_div.sv:26:5
	reg [CNTRW - 1:0] cntr;
	// Trace: src/VX_serial_div.sv:27:5
	reg busy_r;
	// Trace: src/VX_serial_div.sv:28:5
	genvar _gv_i_8;
	generate
		for (_gv_i_8 = 0; _gv_i_8 < LANES; _gv_i_8 = _gv_i_8 + 1) begin : g_setup
			localparam i = _gv_i_8;
			// Trace: src/VX_serial_div.sv:29:9
			wire negate_numer = is_signed && numer[(i * WIDTHN) + (WIDTHN - 1)];
			// Trace: src/VX_serial_div.sv:30:9
			wire negate_denom = is_signed && denom[(i * WIDTHD) + (WIDTHD - 1)];
			// Trace: src/VX_serial_div.sv:31:9
			assign numer_qual[i * WIDTHN+:WIDTHN] = (negate_numer ? -$signed(numer[i * WIDTHN+:WIDTHN]) : numer[i * WIDTHN+:WIDTHN]);
			// Trace: src/VX_serial_div.sv:32:9
			assign denom_qual[i * WIDTHD+:WIDTHD] = (negate_denom ? -$signed(denom[i * WIDTHD+:WIDTHD]) : denom[i * WIDTHD+:WIDTHD]);
			// Trace: src/VX_serial_div.sv:33:9
			assign sub_result[(WIDTHD >= 0 ? 0 : WIDTHD) + (i * (WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD))+:(WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD)] = working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? ((WIDTHN + MIN_ND) >= WIDTHN ? WIDTHN + MIN_ND : ((WIDTHN + MIN_ND) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1) : (WIDTHN + MIN_ND) - ((WIDTHN + MIN_ND) >= WIDTHN ? WIDTHN + MIN_ND : ((WIDTHN + MIN_ND) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? ((WIDTHN + MIN_ND) >= WIDTHN ? WIDTHN + MIN_ND : ((WIDTHN + MIN_ND) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1) : (WIDTHN + MIN_ND) - ((WIDTHN + MIN_ND) >= WIDTHN ? WIDTHN + MIN_ND : ((WIDTHN + MIN_ND) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1))) + ((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)) - 1)-:((WIDTHN + MIN_ND) >= WIDTHN ? ((WIDTHN + MIN_ND) - WIDTHN) + 1 : (WIDTHN - (WIDTHN + MIN_ND)) + 1)] - denom_r[i * WIDTHD+:WIDTHD];
		end
	endgenerate
	// Trace: src/VX_serial_div.sv:35:5
	function automatic signed [CNTRW - 1:0] sv2v_cast_A86AD_signed;
		input reg signed [CNTRW - 1:0] inp;
		sv2v_cast_A86AD_signed = inp;
	endfunction
	always @(posedge clk) begin
		// Trace: src/VX_serial_div.sv:36:9
		if (reset)
			// Trace: src/VX_serial_div.sv:37:13
			busy_r <= 0;
		else begin
			// Trace: src/VX_serial_div.sv:39:13
			if (strobe)
				// Trace: src/VX_serial_div.sv:40:17
				busy_r <= 1;
			if (busy && (cntr == 0))
				// Trace: src/VX_serial_div.sv:43:17
				busy_r <= 0;
		end
		// Trace: src/VX_serial_div.sv:46:9
		cntr <= cntr - sv2v_cast_A86AD_signed(1);
		if (strobe)
			// Trace: src/VX_serial_div.sv:48:13
			cntr <= sv2v_cast_A86AD_signed(WIDTHN - 1);
	end
	// Trace: src/VX_serial_div.sv:51:5
	genvar _gv_i_9;
	generate
		for (_gv_i_9 = 0; _gv_i_9 < LANES; _gv_i_9 = _gv_i_9 + 1) begin : g_div
			localparam i = _gv_i_9;
			// Trace: src/VX_serial_div.sv:52:9
			always @(posedge clk)
				// Trace: src/VX_serial_div.sv:53:13
				if (strobe) begin
					// Trace: src/VX_serial_div.sv:54:17
					working[((WIDTHN + MIN_ND) >= 0 ? 0 : WIDTHN + MIN_ND) + (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND)))+:((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))] <= {{WIDTHD {1'b0}}, numer_qual[i * WIDTHN+:WIDTHN], 1'b0};
					// Trace: src/VX_serial_div.sv:55:17
					denom_r[i * WIDTHD+:WIDTHD] <= denom_qual[i * WIDTHD+:WIDTHD];
					// Trace: src/VX_serial_div.sv:56:17
					inv_quot[i] <= ((denom[i * WIDTHD+:WIDTHD] != 0) && is_signed) && (numer[(i * WIDTHN) + 31] ^ denom[(i * WIDTHD) + 31]);
					// Trace: src/VX_serial_div.sv:57:17
					inv_rem[i] <= is_signed && numer[(i * WIDTHN) + 31];
				end
				else if (busy_r)
					// Trace: src/VX_serial_div.sv:59:17
					working[((WIDTHN + MIN_ND) >= 0 ? 0 : WIDTHN + MIN_ND) + (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND)))+:((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))] <= (sub_result[(i * (WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD)) + (WIDTHD >= 0 ? WIDTHD : WIDTHD - WIDTHD)] ? {working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) - 1 : (WIDTHN + MIN_ND) - ((WIDTHN + MIN_ND) - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) - 1 : (WIDTHN + MIN_ND) - ((WIDTHN + MIN_ND) - 1))) + (WIDTHN + MIN_ND)) - 1)-:WIDTHN + MIN_ND], 1'b0} : {sub_result[(WIDTHD >= 0 ? (i * (WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD)) + (WIDTHD >= 0 ? WIDTHD - 1 : WIDTHD - (WIDTHD - 1)) : (((i * (WIDTHD >= 0 ? WIDTHD + 1 : 1 - WIDTHD)) + (WIDTHD >= 0 ? WIDTHD - 1 : WIDTHD - (WIDTHD - 1))) + WIDTHD) - 1)-:WIDTHD], working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? WIDTHN - 1 : (WIDTHN + MIN_ND) - (WIDTHN - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? WIDTHN - 1 : (WIDTHN + MIN_ND) - (WIDTHN - 1))) + WIDTHN) - 1)-:WIDTHN], 1'b1});
		end
	endgenerate
	// Trace: src/VX_serial_div.sv:64:5
	genvar _gv_i_10;
	generate
		for (_gv_i_10 = 0; _gv_i_10 < LANES; _gv_i_10 = _gv_i_10 + 1) begin : g_output
			localparam i = _gv_i_10;
			// Trace: src/VX_serial_div.sv:65:9
			wire [WIDTHQ - 1:0] q = working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? WIDTHQ - 1 : (WIDTHN + MIN_ND) - (WIDTHQ - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? WIDTHQ - 1 : (WIDTHN + MIN_ND) - (WIDTHQ - 1))) + WIDTHQ) - 1)-:WIDTHQ];
			// Trace: src/VX_serial_div.sv:66:9
			wire [WIDTHR - 1:0] r = working[((WIDTHN + MIN_ND) >= 0 ? (i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? WIDTHN + WIDTHR : ((WIDTHN + WIDTHR) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1) : (WIDTHN + MIN_ND) - ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? WIDTHN + WIDTHR : ((WIDTHN + WIDTHR) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1)) : (((i * ((WIDTHN + MIN_ND) >= 0 ? (WIDTHN + MIN_ND) + 1 : 1 - (WIDTHN + MIN_ND))) + ((WIDTHN + MIN_ND) >= 0 ? ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? WIDTHN + WIDTHR : ((WIDTHN + WIDTHR) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1) : (WIDTHN + MIN_ND) - ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? WIDTHN + WIDTHR : ((WIDTHN + WIDTHR) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1))) + ((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)) - 1)-:((WIDTHN + WIDTHR) >= (WIDTHN + 1) ? ((WIDTHN + WIDTHR) - (WIDTHN + 1)) + 1 : ((WIDTHN + 1) - (WIDTHN + WIDTHR)) + 1)];
			// Trace: src/VX_serial_div.sv:67:9
			assign quotient[i * WIDTHQ+:WIDTHQ] = (inv_quot[i] ? -$signed(q) : q);
			// Trace: src/VX_serial_div.sv:68:9
			assign remainder[i * WIDTHR+:WIDTHR] = (inv_rem[i] ? -$signed(r) : r);
		end
	endgenerate
	// Trace: src/VX_serial_div.sv:70:5
	assign busy = busy_r;
endmodule
module VX_index_buffer (
	clk,
	reset,
	write_addr,
	write_data,
	acquire_en,
	read_addr,
	read_data,
	release_en,
	empty,
	full
);
	// Trace: src/VX_index_buffer.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_index_buffer.sv:3:15
	parameter SIZE = 1;
	// Trace: src/VX_index_buffer.sv:4:15
	parameter LUTRAM = 0;
	// Trace: src/VX_index_buffer.sv:5:15
	parameter ADDRW = (SIZE > 1 ? $clog2(SIZE) : 1);
	// Trace: src/VX_index_buffer.sv:7:5
	input wire clk;
	// Trace: src/VX_index_buffer.sv:8:5
	input wire reset;
	// Trace: src/VX_index_buffer.sv:9:5
	output wire [ADDRW - 1:0] write_addr;
	// Trace: src/VX_index_buffer.sv:10:5
	input wire [DATAW - 1:0] write_data;
	// Trace: src/VX_index_buffer.sv:11:5
	input wire acquire_en;
	// Trace: src/VX_index_buffer.sv:12:5
	input wire [ADDRW - 1:0] read_addr;
	// Trace: src/VX_index_buffer.sv:13:5
	output wire [DATAW - 1:0] read_data;
	// Trace: src/VX_index_buffer.sv:14:5
	input wire release_en;
	// Trace: src/VX_index_buffer.sv:15:5
	output wire empty;
	// Trace: src/VX_index_buffer.sv:16:5
	output wire full;
	// Trace: src/VX_index_buffer.sv:18:5
	VX_allocator #(.SIZE(SIZE)) allocator(
		.clk(clk),
		.reset(reset),
		.acquire_en(acquire_en),
		.acquire_addr(write_addr),
		.release_en(release_en),
		.release_addr(read_addr),
		.empty(empty),
		.full(full)
	);
	// Trace: src/VX_index_buffer.sv:30:5
	VX_dp_ram #(
		.DATAW(DATAW),
		.SIZE(SIZE),
		.LUTRAM(LUTRAM),
		.RDW_MODE("W")
	) data_table(
		.clk(clk),
		.reset(reset),
		.read(1'b1),
		.write(acquire_en),
		.wren(1'b1),
		.waddr(write_addr),
		.wdata(write_data),
		.raddr(read_addr),
		.rdata(read_data)
	);
endmodule
module VX_reduce_tree (
	data_in,
	data_out
);
	// Trace: src/VX_reduce_tree.sv:2:15
	parameter DATAW_IN = 1;
	// Trace: src/VX_reduce_tree.sv:3:15
	parameter DATAW_OUT = DATAW_IN;
	// Trace: src/VX_reduce_tree.sv:4:15
	parameter N = 1;
	// Trace: src/VX_reduce_tree.sv:5:15
	parameter OP = "+";
	// Trace: src/VX_reduce_tree.sv:7:5
	input wire [(N * DATAW_IN) - 1:0] data_in;
	// Trace: src/VX_reduce_tree.sv:8:5
	output wire [DATAW_OUT - 1:0] data_out;
	// Trace: src/VX_reduce_tree.sv:10:5
	function automatic [DATAW_OUT - 1:0] sv2v_cast_0EBAF;
		input reg [DATAW_OUT - 1:0] inp;
		sv2v_cast_0EBAF = inp;
	endfunction
	generate
		if (N == 1) begin : g_passthru
			// Trace: src/VX_reduce_tree.sv:11:9
			assign data_out = sv2v_cast_0EBAF(data_in[0+:DATAW_IN]);
		end
		else begin : g_reduce
			// Trace: src/VX_reduce_tree.sv:13:9
			localparam signed [31:0] N_A = N / 2;
			// Trace: src/VX_reduce_tree.sv:14:9
			localparam signed [31:0] N_B = N - N_A;
			// Trace: src/VX_reduce_tree.sv:15:9
			wire [(N_A * DATAW_IN) - 1:0] in_A;
			// Trace: src/VX_reduce_tree.sv:16:9
			wire [(N_B * DATAW_IN) - 1:0] in_B;
			// Trace: src/VX_reduce_tree.sv:17:9
			wire [DATAW_OUT - 1:0] out_A;
			wire [DATAW_OUT - 1:0] out_B;
			genvar _gv_i_21;
			for (_gv_i_21 = 0; _gv_i_21 < N_A; _gv_i_21 = _gv_i_21 + 1) begin : g_in_A
				localparam i = _gv_i_21;
				// Trace: src/VX_reduce_tree.sv:19:13
				assign in_A[i * DATAW_IN+:DATAW_IN] = data_in[i * DATAW_IN+:DATAW_IN];
			end
			genvar _gv_i_22;
			for (_gv_i_22 = 0; _gv_i_22 < N_B; _gv_i_22 = _gv_i_22 + 1) begin : g_in_B
				localparam i = _gv_i_22;
				// Trace: src/VX_reduce_tree.sv:22:13
				assign in_B[i * DATAW_IN+:DATAW_IN] = data_in[(N_A + i) * DATAW_IN+:DATAW_IN];
			end
			// Trace: src/VX_reduce_tree.sv:24:9
			VX_reduce_tree #(
				.DATAW_IN(DATAW_IN),
				.DATAW_OUT(DATAW_OUT),
				.N(N_A),
				.OP(OP)
			) reduce_A(
				.data_in(in_A),
				.data_out(out_A)
			);
			// Trace: src/VX_reduce_tree.sv:33:9
			VX_reduce_tree #(
				.DATAW_IN(DATAW_IN),
				.DATAW_OUT(DATAW_OUT),
				.N(N_B),
				.OP(OP)
			) reduce_B(
				.data_in(in_B),
				.data_out(out_B)
			);
			if (OP == "+") begin : g_plus
				// Trace: src/VX_reduce_tree.sv:43:13
				assign data_out = out_A + out_B;
			end
			else if (OP == "^") begin : g_xor
				// Trace: src/VX_reduce_tree.sv:45:13
				assign data_out = out_A ^ out_B;
			end
			else if (OP == "&") begin : g_and
				// Trace: src/VX_reduce_tree.sv:47:13
				assign data_out = out_A & out_B;
			end
			else if (OP == "|") begin : g_or
				// Trace: src/VX_reduce_tree.sv:49:13
				assign data_out = out_A | out_B;
			end
		end
	endgenerate
endmodule
module VX_mux (
	data_in,
	sel_in,
	data_out
);
	// Trace: src/VX_mux.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_mux.sv:3:15
	parameter N = 1;
	// Trace: src/VX_mux.sv:4:15
	parameter LN = (N > 1 ? $clog2(N) : 1);
	// Trace: src/VX_mux.sv:6:5
	input wire [(N * DATAW) - 1:0] data_in;
	// Trace: src/VX_mux.sv:7:5
	input wire [LN - 1:0] sel_in;
	// Trace: src/VX_mux.sv:8:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_mux.sv:10:5
	generate
		if (N > 1) begin : g_mux
			// Trace: src/VX_mux.sv:11:9
			assign data_out = data_in[sel_in * DATAW+:DATAW];
		end
		else begin : g_passthru
			// Trace: src/VX_mux.sv:13:9
			assign data_out = data_in;
		end
	endgenerate
endmodule
module VX_pipe_register (
	clk,
	reset,
	enable,
	data_in,
	data_out
);
	// Trace: src/VX_pipe_register.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_pipe_register.sv:3:15
	parameter RESETW = 0;
	// Trace: src/VX_pipe_register.sv:4:15
	parameter DEPTH = 1;
	// Trace: src/VX_pipe_register.sv:5:15
	parameter [(RESETW > 0 ? RESETW : 1) - 1:0] INIT_VALUE = {(RESETW > 0 ? RESETW : 1) {1'b0}};
	// Trace: src/VX_pipe_register.sv:7:5
	input wire clk;
	// Trace: src/VX_pipe_register.sv:8:5
	input wire reset;
	// Trace: src/VX_pipe_register.sv:9:5
	input wire enable;
	// Trace: src/VX_pipe_register.sv:10:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_pipe_register.sv:11:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_pipe_register.sv:13:5
	VX_shift_register #(
		.DATAW(DATAW),
		.RESETW(RESETW),
		.DEPTH(DEPTH),
		.INIT_VALUE(INIT_VALUE)
	) g_shift_register(
		.clk(clk),
		.reset(reset),
		.enable(enable),
		.data_in(data_in),
		.data_out(data_out)
	);
endmodule
// removed module with interface ports: VX_alu_unit
// removed module with interface ports: VX_lsu_mem_arb
module VX_stream_pack (
	clk,
	reset,
	valid_in,
	data_in,
	tag_in,
	ready_in,
	valid_out,
	mask_out,
	data_out,
	tag_out,
	ready_out
);
	// Trace: src/VX_stream_pack.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_stream_pack.sv:3:15
	parameter DATA_WIDTH = 1;
	// Trace: src/VX_stream_pack.sv:4:15
	parameter TAG_WIDTH = 1;
	// Trace: src/VX_stream_pack.sv:5:15
	parameter TAG_SEL_BITS = 0;
	// Trace: src/VX_stream_pack.sv:6:15
	parameter ARBITER = "P";
	// Trace: src/VX_stream_pack.sv:7:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_stream_pack.sv:9:5
	input wire clk;
	// Trace: src/VX_stream_pack.sv:10:5
	input wire reset;
	// Trace: src/VX_stream_pack.sv:11:5
	input wire [NUM_REQS - 1:0] valid_in;
	// Trace: src/VX_stream_pack.sv:12:5
	input wire [(NUM_REQS * DATA_WIDTH) - 1:0] data_in;
	// Trace: src/VX_stream_pack.sv:13:5
	input wire [(NUM_REQS * TAG_WIDTH) - 1:0] tag_in;
	// Trace: src/VX_stream_pack.sv:14:5
	output wire [NUM_REQS - 1:0] ready_in;
	// Trace: src/VX_stream_pack.sv:15:5
	output wire valid_out;
	// Trace: src/VX_stream_pack.sv:16:5
	output wire [NUM_REQS - 1:0] mask_out;
	// Trace: src/VX_stream_pack.sv:17:5
	output wire [(NUM_REQS * DATA_WIDTH) - 1:0] data_out;
	// Trace: src/VX_stream_pack.sv:18:5
	output wire [TAG_WIDTH - 1:0] tag_out;
	// Trace: src/VX_stream_pack.sv:19:5
	input wire ready_out;
	// Trace: src/VX_stream_pack.sv:21:5
	generate
		if (NUM_REQS > 1) begin : g_pack
			// Trace: src/VX_stream_pack.sv:22:9
			localparam LOG_NUM_REQS = $clog2(NUM_REQS);
			// Trace: src/VX_stream_pack.sv:23:9
			wire [LOG_NUM_REQS - 1:0] grant_index;
			// Trace: src/VX_stream_pack.sv:24:9
			wire grant_valid;
			// Trace: src/VX_stream_pack.sv:25:9
			wire grant_ready;
			// Trace: src/VX_stream_pack.sv:26:9
			VX_generic_arbiter #(
				.NUM_REQS(NUM_REQS),
				.TYPE(ARBITER)
			) arbiter(
				.clk(clk),
				.reset(reset),
				.requests(valid_in),
				.grant_valid(grant_valid),
				.grant_index(grant_index),
				.grant_onehot(),
				.grant_ready(grant_ready)
			);
			// Trace: src/VX_stream_pack.sv:38:9
			wire [TAG_WIDTH - 1:0] tag_sel = tag_in[grant_index * TAG_WIDTH+:TAG_WIDTH];
			// Trace: src/VX_stream_pack.sv:39:9
			wire [NUM_REQS - 1:0] tag_matches;
			genvar _gv_i_28;
			for (_gv_i_28 = 0; _gv_i_28 < NUM_REQS; _gv_i_28 = _gv_i_28 + 1) begin : g_tag_matches
				localparam i = _gv_i_28;
				// Trace: src/VX_stream_pack.sv:41:13
				assign tag_matches[i] = tag_in[(i * TAG_WIDTH) + (TAG_SEL_BITS - 1)-:TAG_SEL_BITS] == tag_sel[TAG_SEL_BITS - 1:0];
			end
			genvar _gv_i_29;
			for (_gv_i_29 = 0; _gv_i_29 < NUM_REQS; _gv_i_29 = _gv_i_29 + 1) begin : g_ready_in
				localparam i = _gv_i_29;
				// Trace: src/VX_stream_pack.sv:44:13
				assign ready_in[i] = grant_ready & tag_matches[i];
			end
			// Trace: src/VX_stream_pack.sv:46:9
			wire [NUM_REQS - 1:0] mask_sel = valid_in & tag_matches;
			// Trace: src/VX_stream_pack.sv:47:9
			VX_elastic_buffer #(
				.DATAW((NUM_REQS + TAG_WIDTH) + (NUM_REQS * DATA_WIDTH)),
				.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
				.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
			) out_buf(
				.clk(clk),
				.reset(reset),
				.valid_in(grant_valid),
				.data_in({mask_sel, tag_sel, data_in}),
				.ready_in(grant_ready),
				.valid_out(valid_out),
				.data_out({mask_out, tag_out, data_out}),
				.ready_out(ready_out)
			);
		end
		else begin : g_passthru
			// Trace: src/VX_stream_pack.sv:62:9
			assign valid_out = valid_in;
			// Trace: src/VX_stream_pack.sv:63:9
			assign mask_out = 1'b1;
			// Trace: src/VX_stream_pack.sv:64:9
			assign data_out = data_in;
			// Trace: src/VX_stream_pack.sv:65:9
			assign tag_out = tag_in;
			// Trace: src/VX_stream_pack.sv:66:9
			assign ready_in = ready_out;
		end
	endgenerate
endmodule
module VX_allocator (
	clk,
	reset,
	acquire_en,
	acquire_addr,
	release_en,
	release_addr,
	empty,
	full
);
	// Trace: src/VX_allocator.sv:2:15
	parameter SIZE = 1;
	// Trace: src/VX_allocator.sv:3:15
	parameter ADDRW = (SIZE > 1 ? $clog2(SIZE) : 1);
	// Trace: src/VX_allocator.sv:5:5
	input wire clk;
	// Trace: src/VX_allocator.sv:6:5
	input wire reset;
	// Trace: src/VX_allocator.sv:7:5
	input wire acquire_en;
	// Trace: src/VX_allocator.sv:8:5
	output wire [ADDRW - 1:0] acquire_addr;
	// Trace: src/VX_allocator.sv:9:5
	input wire release_en;
	// Trace: src/VX_allocator.sv:10:5
	input wire [ADDRW - 1:0] release_addr;
	// Trace: src/VX_allocator.sv:11:5
	output wire empty;
	// Trace: src/VX_allocator.sv:12:5
	output wire full;
	// Trace: src/VX_allocator.sv:14:5
	reg [SIZE - 1:0] free_slots;
	reg [SIZE - 1:0] free_slots_n;
	// Trace: src/VX_allocator.sv:15:5
	reg [ADDRW - 1:0] acquire_addr_r;
	// Trace: src/VX_allocator.sv:16:5
	reg empty_r;
	reg full_r;
	// Trace: src/VX_allocator.sv:17:5
	wire [ADDRW - 1:0] free_index;
	// Trace: src/VX_allocator.sv:18:5
	wire free_valid;
	// Trace: src/VX_allocator.sv:19:5
	always @(*) begin
		// Trace: src/VX_allocator.sv:20:9
		free_slots_n = free_slots;
		// Trace: src/VX_allocator.sv:21:9
		if (release_en)
			// Trace: src/VX_allocator.sv:22:13
			free_slots_n[release_addr] = 1;
		if (acquire_en)
			// Trace: src/VX_allocator.sv:25:13
			free_slots_n[acquire_addr_r] = 0;
	end
	// Trace: src/VX_allocator.sv:28:5
	VX_priority_encoder #(.N(SIZE)) free_slots_sel(
		.data_in(free_slots_n),
		.index_out(free_index),
		.valid_out(free_valid),
		.onehot_out()
	);
	// Trace: src/VX_allocator.sv:36:5
	function automatic [ADDRW - 1:0] sv2v_cast_8BB5D;
		input reg [ADDRW - 1:0] inp;
		sv2v_cast_8BB5D = inp;
	endfunction
	always @(posedge clk)
		// Trace: src/VX_allocator.sv:37:9
		if (reset) begin
			// Trace: src/VX_allocator.sv:38:13
			acquire_addr_r <= sv2v_cast_8BB5D(1'b0);
			// Trace: src/VX_allocator.sv:39:13
			free_slots <= {SIZE {1'b1}};
			// Trace: src/VX_allocator.sv:40:13
			empty_r <= 1'b1;
			// Trace: src/VX_allocator.sv:41:13
			full_r <= 1'b0;
		end
		else begin
			// Trace: src/VX_allocator.sv:43:13
			if (release_en)
				;
			if (acquire_en)
				;
			if (acquire_en || (release_en && full_r))
				// Trace: src/VX_allocator.sv:50:17
				acquire_addr_r <= free_index;
			// Trace: src/VX_allocator.sv:52:13
			free_slots <= free_slots_n;
			// Trace: src/VX_allocator.sv:53:13
			empty_r <= &free_slots_n;
			// Trace: src/VX_allocator.sv:54:13
			full_r <= ~free_valid;
		end
	// Trace: src/VX_allocator.sv:57:5
	assign acquire_addr = acquire_addr_r;
	// Trace: src/VX_allocator.sv:58:5
	assign empty = empty_r;
	// Trace: src/VX_allocator.sv:59:5
	assign full = full_r;
endmodule
// removed interface: VX_commit_sched_if
module VX_bits_insert (
	data_in,
	ins_in,
	data_out
);
	// Trace: src/VX_bits_insert.sv:2:15
	parameter N = 1;
	// Trace: src/VX_bits_insert.sv:3:15
	parameter S = 1;
	// Trace: src/VX_bits_insert.sv:4:15
	parameter POS = 0;
	// Trace: src/VX_bits_insert.sv:6:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_bits_insert.sv:7:5
	input wire [(S > 0 ? S : 1) - 1:0] ins_in;
	// Trace: src/VX_bits_insert.sv:8:5
	output wire [(N + S) - 1:0] data_out;
	// Trace: src/VX_bits_insert.sv:10:5
	generate
		if (S == 0) begin : g_passthru
			// Trace: src/VX_bits_insert.sv:11:9
			assign data_out = data_in;
		end
		else begin : g_insert
			if (POS == 0) begin : g_pos_0
				// Trace: src/VX_bits_insert.sv:14:13
				assign data_out = {data_in, ins_in};
			end
			else if (POS == N) begin : g_pos_N
				// Trace: src/VX_bits_insert.sv:16:13
				assign data_out = {ins_in, data_in};
			end
			else begin : g_pos
				// Trace: src/VX_bits_insert.sv:18:13
				assign data_out = {data_in[N - 1:POS], ins_in, data_in[POS - 1:0]};
			end
		end
	endgenerate
endmodule
module VX_find_first (
	data_in,
	valid_in,
	data_out,
	valid_out
);
	// Trace: src/VX_find_first.sv:2:15
	parameter N = 1;
	// Trace: src/VX_find_first.sv:3:15
	parameter DATAW = 1;
	// Trace: src/VX_find_first.sv:4:15
	parameter REVERSE = 0;
	// Trace: src/VX_find_first.sv:6:5
	input wire [(N * DATAW) - 1:0] data_in;
	// Trace: src/VX_find_first.sv:7:5
	input wire [N - 1:0] valid_in;
	// Trace: src/VX_find_first.sv:8:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_find_first.sv:9:5
	output wire valid_out;
	// Trace: src/VX_find_first.sv:11:5
	localparam LOGN = $clog2(N);
	// Trace: src/VX_find_first.sv:12:5
	localparam TL = (1 << LOGN) - 1;
	// Trace: src/VX_find_first.sv:13:5
	localparam TN = (1 << (LOGN + 1)) - 1;
	// Trace: src/VX_find_first.sv:14:5
	wire s_n [0:TN - 1];
	// Trace: src/VX_find_first.sv:15:5
	wire [DATAW - 1:0] d_n [0:TN - 1];
	// Trace: src/VX_find_first.sv:16:5
	genvar _gv_i_32;
	generate
		for (_gv_i_32 = 0; _gv_i_32 < N; _gv_i_32 = _gv_i_32 + 1) begin : g_fill
			localparam i = _gv_i_32;
			// Trace: src/VX_find_first.sv:17:9
			assign s_n[TL + i] = (REVERSE ? valid_in[(N - 1) - i] : valid_in[i]);
			// Trace: src/VX_find_first.sv:18:9
			assign d_n[TL + i] = (REVERSE ? data_in[((N - 1) - i) * DATAW+:DATAW] : data_in[i * DATAW+:DATAW]);
		end
	endgenerate
	// Trace: src/VX_find_first.sv:20:5
	generate
		if (TL < (TN - N)) begin : g_padding
			genvar _gv_i_33;
			for (_gv_i_33 = TL + N; _gv_i_33 < TN; _gv_i_33 = _gv_i_33 + 1) begin : g_i
				localparam i = _gv_i_33;
				// Trace: src/VX_find_first.sv:22:13
				assign s_n[i] = 0;
				// Trace: src/VX_find_first.sv:23:13
				assign d_n[i] = 1'sb0;
			end
		end
	endgenerate
	// Trace: src/VX_find_first.sv:26:5
	genvar _gv_j_2;
	generate
		for (_gv_j_2 = 0; _gv_j_2 < LOGN; _gv_j_2 = _gv_j_2 + 1) begin : g_scan
			localparam j = _gv_j_2;
			// Trace: src/VX_find_first.sv:27:9
			localparam I = 1 << j;
			genvar _gv_i_34;
			for (_gv_i_34 = 0; _gv_i_34 < I; _gv_i_34 = _gv_i_34 + 1) begin : g_i
				localparam i = _gv_i_34;
				// Trace: src/VX_find_first.sv:29:13
				localparam K = (I + i) - 1;
				// Trace: src/VX_find_first.sv:30:13
				assign s_n[K] = s_n[(2 * K) + 2] | s_n[(2 * K) + 1];
				// Trace: src/VX_find_first.sv:31:13
				assign d_n[K] = (s_n[(2 * K) + 1] ? d_n[(2 * K) + 1] : d_n[(2 * K) + 2]);
			end
		end
	endgenerate
	// Trace: src/VX_find_first.sv:34:5
	assign valid_out = s_n[0];
	// Trace: src/VX_find_first.sv:35:5
	assign data_out = d_n[0];
endmodule
// removed module with interface ports: VX_dispatch_unit
// removed interface: VX_gbar_bus_if
// removed module with interface ports: VX_cache_wrap
module VX_pipe_buffer (
	clk,
	reset,
	valid_in,
	ready_in,
	data_in,
	data_out,
	ready_out,
	valid_out
);
	// Trace: src/VX_pipe_buffer.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_pipe_buffer.sv:3:15
	parameter RESETW = 0;
	// Trace: src/VX_pipe_buffer.sv:4:15
	parameter DEPTH = 1;
	// Trace: src/VX_pipe_buffer.sv:6:5
	input wire clk;
	// Trace: src/VX_pipe_buffer.sv:7:5
	input wire reset;
	// Trace: src/VX_pipe_buffer.sv:8:5
	input wire valid_in;
	// Trace: src/VX_pipe_buffer.sv:9:5
	output wire ready_in;
	// Trace: src/VX_pipe_buffer.sv:10:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_pipe_buffer.sv:11:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_pipe_buffer.sv:12:5
	input wire ready_out;
	// Trace: src/VX_pipe_buffer.sv:13:5
	output wire valid_out;
	// Trace: src/VX_pipe_buffer.sv:15:5
	generate
		if (DEPTH == 0) begin : g_passthru
			// Trace: src/VX_pipe_buffer.sv:16:9
			assign ready_in = ready_out;
			// Trace: src/VX_pipe_buffer.sv:17:9
			assign valid_out = valid_in;
			// Trace: src/VX_pipe_buffer.sv:18:9
			assign data_out = data_in;
		end
		else begin : g_register
			// Trace: src/VX_pipe_buffer.sv:20:9
			wire [DEPTH:0] valid;
			// Trace: src/VX_pipe_buffer.sv:21:9
			wire ready [0:DEPTH + 0];
			// Trace: src/VX_pipe_buffer.sv:22:9
			wire [(DEPTH >= 0 ? ((DEPTH + 1) * DATAW) - 1 : ((1 - DEPTH) * DATAW) + ((DEPTH * DATAW) - 1)):(DEPTH >= 0 ? 0 : DEPTH * DATAW)] data;
			// Trace: src/VX_pipe_buffer.sv:23:9
			assign valid[0] = valid_in;
			// Trace: src/VX_pipe_buffer.sv:24:9
			assign data[(DEPTH >= 0 ? 0 : DEPTH) * DATAW+:DATAW] = data_in;
			// Trace: src/VX_pipe_buffer.sv:25:9
			assign ready_in = ready[0];
			genvar _gv_i_47;
			for (_gv_i_47 = 0; _gv_i_47 < DEPTH; _gv_i_47 = _gv_i_47 + 1) begin : g_pipe_regs
				localparam i = _gv_i_47;
				// Trace: src/VX_pipe_buffer.sv:27:13
				assign ready[i] = ready[i + 1] || ~valid[i + 1];
				// Trace: src/VX_pipe_buffer.sv:28:13
				VX_pipe_register #(
					.DATAW(1 + DATAW),
					.RESETW(1 + RESETW)
				) pipe_register(
					.clk(clk),
					.reset(reset),
					.enable(ready[i]),
					.data_in({valid[i], data[(DEPTH >= 0 ? i : DEPTH - i) * DATAW+:DATAW]}),
					.data_out({valid[i + 1], data[(DEPTH >= 0 ? i + 1 : DEPTH - (i + 1)) * DATAW+:DATAW]})
				);
			end
			// Trace: src/VX_pipe_buffer.sv:39:9
			assign valid_out = valid[DEPTH];
			// Trace: src/VX_pipe_buffer.sv:40:9
			assign data_out = data[(DEPTH >= 0 ? DEPTH : DEPTH - DEPTH) * DATAW+:DATAW];
			// Trace: src/VX_pipe_buffer.sv:41:9
			assign ready[DEPTH] = ready_out;
		end
	endgenerate
endmodule
module VX_bits_remove (
	data_in,
	sel_out,
	data_out
);
	// Trace: src/VX_bits_remove.sv:2:15
	parameter N = 2;
	// Trace: src/VX_bits_remove.sv:3:15
	parameter S = 1;
	// Trace: src/VX_bits_remove.sv:4:15
	parameter POS = 0;
	// Trace: src/VX_bits_remove.sv:6:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_bits_remove.sv:7:5
	output wire [(S > 0 ? S : 1) - 1:0] sel_out;
	// Trace: src/VX_bits_remove.sv:8:5
	output wire [(N - S) - 1:0] data_out;
	// Trace: src/VX_bits_remove.sv:10:5
	generate
		if (S == 0) begin : g_passthru
			// Trace: src/VX_bits_remove.sv:11:9
			assign sel_out = 0;
			// Trace: src/VX_bits_remove.sv:12:9
			assign data_out = data_in;
		end
		else if (POS == 0) begin : g_pos_0
			// Trace: src/VX_bits_remove.sv:14:9
			assign sel_out = data_in[0+:S];
			// Trace: src/VX_bits_remove.sv:15:9
			assign data_out = data_in[N - 1:S];
		end
		else if ((POS + S) == N) begin : g_pos_N
			// Trace: src/VX_bits_remove.sv:17:9
			assign sel_out = data_in[POS+:S];
			// Trace: src/VX_bits_remove.sv:18:9
			assign data_out = data_in[POS - 1:0];
		end
		else begin : g_pos
			// Trace: src/VX_bits_remove.sv:20:9
			assign sel_out = data_in[POS+:S];
			// Trace: src/VX_bits_remove.sv:21:9
			assign data_out = {data_in[N - 1:POS + S], data_in[POS - 1:0]};
		end
	endgenerate
endmodule
// removed interface: VX_ibuffer_if
// removed module with interface ports: VX_lmem_switch
// removed module with interface ports: VX_issue
module VX_priority_encoder (
	data_in,
	onehot_out,
	index_out,
	valid_out
);
	// Trace: src/VX_priority_encoder.sv:2:15
	parameter N = 1;
	// Trace: src/VX_priority_encoder.sv:3:15
	parameter REVERSE = 0;
	// Trace: src/VX_priority_encoder.sv:4:15
	parameter MODEL = 1;
	// Trace: src/VX_priority_encoder.sv:5:15
	parameter LN = (N > 1 ? $clog2(N) : 1);
	// Trace: src/VX_priority_encoder.sv:7:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_priority_encoder.sv:8:5
	output wire [N - 1:0] onehot_out;
	// Trace: src/VX_priority_encoder.sv:9:5
	output wire [LN - 1:0] index_out;
	// Trace: src/VX_priority_encoder.sv:10:5
	output wire valid_out;
	// Trace: src/VX_priority_encoder.sv:12:5
	function automatic signed [LN - 1:0] sv2v_cast_83428_signed;
		input reg signed [LN - 1:0] inp;
		sv2v_cast_83428_signed = inp;
	endfunction
	function automatic signed [N - 1:0] sv2v_cast_AC047_signed;
		input reg signed [N - 1:0] inp;
		sv2v_cast_AC047_signed = inp;
	endfunction
	generate
		if (REVERSE) begin : g_msb
			if (N == 1) begin : g_n1
				// Trace: src/VX_priority_encoder.sv:14:13
				assign onehot_out = data_in;
				// Trace: src/VX_priority_encoder.sv:15:13
				assign index_out = 1'sb0;
				// Trace: src/VX_priority_encoder.sv:16:13
				assign valid_out = data_in;
			end
			else if (N == 2) begin : g_n2
				// Trace: src/VX_priority_encoder.sv:18:13
				assign onehot_out = {data_in[1], data_in[0] & ~data_in[1]};
				// Trace: src/VX_priority_encoder.sv:19:13
				assign index_out = data_in[1];
				// Trace: src/VX_priority_encoder.sv:20:13
				assign valid_out = |data_in;
			end
			else if (MODEL != 0) begin : g_model1
				// Trace: src/VX_priority_encoder.sv:22:13
				wire [N - 1:0] higher_pri_regs;
				// Trace: src/VX_priority_encoder.sv:23:13
				assign higher_pri_regs[N - 1] = 1'b0;
				genvar _gv_i_49;
				for (_gv_i_49 = N - 2; _gv_i_49 >= 0; _gv_i_49 = _gv_i_49 - 1) begin : g_higher_pri_regs
					localparam i = _gv_i_49;
					// Trace: src/VX_priority_encoder.sv:25:17
					assign higher_pri_regs[i] = higher_pri_regs[i + 1] | data_in[i + 1];
				end
				// Trace: src/VX_priority_encoder.sv:27:13
				assign onehot_out = data_in & ~higher_pri_regs;
				// Trace: src/VX_priority_encoder.sv:28:13
				wire [(N * LN) - 1:0] indices;
				genvar _gv_i_50;
				for (_gv_i_50 = 0; _gv_i_50 < N; _gv_i_50 = _gv_i_50 + 1) begin : g_indices
					localparam i = _gv_i_50;
					// Trace: src/VX_priority_encoder.sv:30:17
					assign indices[i * LN+:LN] = sv2v_cast_83428_signed(i);
				end
				// Trace: src/VX_priority_encoder.sv:32:13
				VX_find_first #(
					.N(N),
					.DATAW(LN),
					.REVERSE(1)
				) find_first(
					.valid_in(data_in),
					.data_in(indices),
					.data_out(index_out),
					.valid_out(valid_out)
				);
			end
			else begin : g_model0
				// Trace: src/VX_priority_encoder.sv:43:13
				reg [LN - 1:0] index_w;
				// Trace: src/VX_priority_encoder.sv:44:13
				reg [N - 1:0] onehot_w;
				// Trace: src/VX_priority_encoder.sv:45:13
				always @(*) begin
					// Trace: src/VX_priority_encoder.sv:46:17
					index_w = 1'sbx;
					// Trace: src/VX_priority_encoder.sv:47:17
					onehot_w = 1'sbx;
					// Trace: src/VX_priority_encoder.sv:48:17
					begin : sv2v_autoblock_1
						// Trace: src/VX_priority_encoder.sv:48:22
						integer i;
						// Trace: src/VX_priority_encoder.sv:48:22
						for (i = 0; i < (N - 1); i = i + 1)
							begin
								// Trace: src/VX_priority_encoder.sv:49:21
								if (data_in[i]) begin
									// Trace: src/VX_priority_encoder.sv:50:25
									index_w = sv2v_cast_83428_signed(i);
									// Trace: src/VX_priority_encoder.sv:51:25
									onehot_w = sv2v_cast_AC047_signed(1) << i;
								end
							end
					end
				end
				// Trace: src/VX_priority_encoder.sv:55:13
				assign index_out = index_w;
				// Trace: src/VX_priority_encoder.sv:56:13
				assign onehot_out = onehot_w;
				// Trace: src/VX_priority_encoder.sv:57:13
				assign valid_out = |data_in;
			end
		end
		else begin : g_lsb
			if (N == 1) begin : g_n1
				// Trace: src/VX_priority_encoder.sv:61:13
				assign onehot_out = data_in;
				// Trace: src/VX_priority_encoder.sv:62:13
				assign index_out = 1'sb0;
				// Trace: src/VX_priority_encoder.sv:63:13
				assign valid_out = data_in;
			end
			else if (N == 2) begin : g_n2
				// Trace: src/VX_priority_encoder.sv:65:13
				assign onehot_out = {data_in[1] && ~data_in[0], data_in[0]};
				// Trace: src/VX_priority_encoder.sv:66:13
				assign index_out = ~data_in[0];
				// Trace: src/VX_priority_encoder.sv:67:13
				assign valid_out = |data_in;
			end
			else if (MODEL == 1) begin : g_model1
				// Trace: src/VX_priority_encoder.sv:69:13
				wire [N - 1:0] higher_pri_regs;
				// Trace: src/VX_priority_encoder.sv:70:13
				assign higher_pri_regs[0] = 1'b0;
				genvar _gv_i_51;
				for (_gv_i_51 = 1; _gv_i_51 < N; _gv_i_51 = _gv_i_51 + 1) begin : g_higher_pri_regs
					localparam i = _gv_i_51;
					// Trace: src/VX_priority_encoder.sv:72:17
					assign higher_pri_regs[i] = higher_pri_regs[i - 1] | data_in[i - 1];
				end
				// Trace: src/VX_priority_encoder.sv:74:13
				assign onehot_out[N - 1:0] = data_in[N - 1:0] & ~higher_pri_regs[N - 1:0];
				// Trace: src/VX_priority_encoder.sv:75:13
				VX_lzc #(
					.N(N),
					.REVERSE(1)
				) lzc(
					.data_in(data_in),
					.data_out(index_out),
					.valid_out(valid_out)
				);
			end
			else if (MODEL == 2) begin : g_model2
				// Trace: src/VX_priority_encoder.sv:84:13
				wire [N - 1:0] scan_lo;
				// Trace: src/VX_priority_encoder.sv:85:13
				VX_scan #(
					.N(N),
					.OP("|")
				) scan(
					.data_in(data_in),
					.data_out(scan_lo)
				);
				// Trace: src/VX_priority_encoder.sv:92:13
				assign onehot_out = scan_lo & {~scan_lo[N - 2:0], 1'b1};
				// Trace: src/VX_priority_encoder.sv:93:13
				VX_lzc #(
					.N(N),
					.REVERSE(1)
				) lzc(
					.data_in(data_in),
					.data_out(index_out),
					.valid_out(valid_out)
				);
			end
			else if (MODEL == 3) begin : g_model3
				// Trace: src/VX_priority_encoder.sv:102:13
				assign onehot_out = data_in & -data_in;
				// Trace: src/VX_priority_encoder.sv:103:13
				VX_lzc #(
					.N(N),
					.REVERSE(1)
				) lzc(
					.data_in(data_in),
					.data_out(index_out),
					.valid_out(valid_out)
				);
			end
			else begin : g_model0
				// Trace: src/VX_priority_encoder.sv:112:13
				reg [LN - 1:0] index_w;
				// Trace: src/VX_priority_encoder.sv:113:13
				reg [N - 1:0] onehot_w;
				// Trace: src/VX_priority_encoder.sv:114:13
				always @(*) begin
					// Trace: src/VX_priority_encoder.sv:115:17
					index_w = 1'sbx;
					// Trace: src/VX_priority_encoder.sv:116:17
					onehot_w = 1'sbx;
					// Trace: src/VX_priority_encoder.sv:117:17
					begin : sv2v_autoblock_2
						// Trace: src/VX_priority_encoder.sv:117:22
						integer i;
						// Trace: src/VX_priority_encoder.sv:117:22
						for (i = N - 1; i >= 0; i = i - 1)
							begin
								// Trace: src/VX_priority_encoder.sv:118:21
								if (data_in[i]) begin
									// Trace: src/VX_priority_encoder.sv:119:25
									index_w = sv2v_cast_83428_signed(i);
									// Trace: src/VX_priority_encoder.sv:120:25
									onehot_w = sv2v_cast_AC047_signed(1) << i;
								end
							end
					end
				end
				// Trace: src/VX_priority_encoder.sv:124:13
				assign index_out = index_w;
				// Trace: src/VX_priority_encoder.sv:125:13
				assign onehot_out = onehot_w;
				// Trace: src/VX_priority_encoder.sv:126:13
				assign valid_out = |data_in;
			end
		end
	endgenerate
endmodule
module VX_mem_scheduler (
	clk,
	reset,
	core_req_valid,
	core_req_rw,
	core_req_mask,
	core_req_byteen,
	core_req_addr,
	core_req_flags,
	core_req_data,
	core_req_tag,
	core_req_ready,
	req_queue_empty,
	req_queue_rw_notify,
	core_rsp_valid,
	core_rsp_mask,
	core_rsp_data,
	core_rsp_tag,
	core_rsp_sop,
	core_rsp_eop,
	core_rsp_ready,
	mem_req_valid,
	mem_req_rw,
	mem_req_mask,
	mem_req_byteen,
	mem_req_addr,
	mem_req_flags,
	mem_req_data,
	mem_req_tag,
	mem_req_ready,
	mem_rsp_valid,
	mem_rsp_mask,
	mem_rsp_data,
	mem_rsp_tag,
	mem_rsp_ready
);
	// Trace: src/VX_mem_scheduler.sv:2:15
	parameter INSTANCE_ID = "";
	// Trace: src/VX_mem_scheduler.sv:3:15
	parameter CORE_REQS = 1;
	// Trace: src/VX_mem_scheduler.sv:4:15
	parameter MEM_CHANNELS = 1;
	// Trace: src/VX_mem_scheduler.sv:5:15
	parameter WORD_SIZE = 4;
	// Trace: src/VX_mem_scheduler.sv:6:15
	parameter LINE_SIZE = WORD_SIZE;
	// Trace: src/VX_mem_scheduler.sv:7:15
	parameter ADDR_WIDTH = 32 - $clog2(WORD_SIZE);
	// Trace: src/VX_mem_scheduler.sv:8:15
	parameter FLAGS_WIDTH = 0;
	// Trace: src/VX_mem_scheduler.sv:9:15
	parameter TAG_WIDTH = 8;
	// Trace: src/VX_mem_scheduler.sv:10:15
	parameter UUID_WIDTH = 0;
	// Trace: src/VX_mem_scheduler.sv:11:15
	parameter CORE_QUEUE_SIZE = 8;
	// Trace: src/VX_mem_scheduler.sv:12:15
	parameter MEM_QUEUE_SIZE = CORE_QUEUE_SIZE;
	// Trace: src/VX_mem_scheduler.sv:13:15
	parameter RSP_PARTIAL = 0;
	// Trace: src/VX_mem_scheduler.sv:14:15
	parameter CORE_OUT_BUF = 0;
	// Trace: src/VX_mem_scheduler.sv:15:15
	parameter MEM_OUT_BUF = 0;
	// Trace: src/VX_mem_scheduler.sv:16:15
	parameter WORD_WIDTH = WORD_SIZE * 8;
	// Trace: src/VX_mem_scheduler.sv:17:15
	parameter LINE_WIDTH = LINE_SIZE * 8;
	// Trace: src/VX_mem_scheduler.sv:18:15
	parameter COALESCE_ENABLE = (CORE_REQS > 1) && (LINE_SIZE != WORD_SIZE);
	// Trace: src/VX_mem_scheduler.sv:19:15
	parameter PER_LINE_REQS = LINE_SIZE / WORD_SIZE;
	// Trace: src/VX_mem_scheduler.sv:20:15
	parameter MERGED_REQS = CORE_REQS / PER_LINE_REQS;
	// Trace: src/VX_mem_scheduler.sv:21:15
	parameter MEM_BATCHES = ((MERGED_REQS + MEM_CHANNELS) - 1) / MEM_CHANNELS;
	// Trace: src/VX_mem_scheduler.sv:22:15
	parameter MEM_BATCH_BITS = $clog2(MEM_BATCHES);
	// Trace: src/VX_mem_scheduler.sv:23:15
	parameter MEM_QUEUE_ADDRW = $clog2((COALESCE_ENABLE ? MEM_QUEUE_SIZE : CORE_QUEUE_SIZE));
	// Trace: src/VX_mem_scheduler.sv:24:15
	parameter MEM_ADDR_WIDTH = ADDR_WIDTH - $clog2(PER_LINE_REQS);
	// Trace: src/VX_mem_scheduler.sv:25:15
	parameter MEM_TAG_WIDTH = (UUID_WIDTH + MEM_QUEUE_ADDRW) + MEM_BATCH_BITS;
	// Trace: src/VX_mem_scheduler.sv:26:15
	parameter CORE_QUEUE_ADDRW = $clog2(CORE_QUEUE_SIZE);
	// Trace: src/VX_mem_scheduler.sv:28:5
	input wire clk;
	// Trace: src/VX_mem_scheduler.sv:29:5
	input wire reset;
	// Trace: src/VX_mem_scheduler.sv:30:5
	input wire core_req_valid;
	// Trace: src/VX_mem_scheduler.sv:31:5
	input wire core_req_rw;
	// Trace: src/VX_mem_scheduler.sv:32:5
	input wire [CORE_REQS - 1:0] core_req_mask;
	// Trace: src/VX_mem_scheduler.sv:33:5
	input wire [(CORE_REQS * WORD_SIZE) - 1:0] core_req_byteen;
	// Trace: src/VX_mem_scheduler.sv:34:5
	input wire [(CORE_REQS * ADDR_WIDTH) - 1:0] core_req_addr;
	// Trace: src/VX_mem_scheduler.sv:35:5
	input wire [(CORE_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] core_req_flags;
	// Trace: src/VX_mem_scheduler.sv:36:5
	input wire [(CORE_REQS * WORD_WIDTH) - 1:0] core_req_data;
	// Trace: src/VX_mem_scheduler.sv:37:5
	input wire [TAG_WIDTH - 1:0] core_req_tag;
	// Trace: src/VX_mem_scheduler.sv:38:5
	output wire core_req_ready;
	// Trace: src/VX_mem_scheduler.sv:39:5
	output wire req_queue_empty;
	// Trace: src/VX_mem_scheduler.sv:40:5
	output wire req_queue_rw_notify;
	// Trace: src/VX_mem_scheduler.sv:41:5
	output wire core_rsp_valid;
	// Trace: src/VX_mem_scheduler.sv:42:5
	output wire [CORE_REQS - 1:0] core_rsp_mask;
	// Trace: src/VX_mem_scheduler.sv:43:5
	output wire [(CORE_REQS * WORD_WIDTH) - 1:0] core_rsp_data;
	// Trace: src/VX_mem_scheduler.sv:44:5
	output wire [TAG_WIDTH - 1:0] core_rsp_tag;
	// Trace: src/VX_mem_scheduler.sv:45:5
	output wire core_rsp_sop;
	// Trace: src/VX_mem_scheduler.sv:46:5
	output wire core_rsp_eop;
	// Trace: src/VX_mem_scheduler.sv:47:5
	input wire core_rsp_ready;
	// Trace: src/VX_mem_scheduler.sv:48:5
	output wire mem_req_valid;
	// Trace: src/VX_mem_scheduler.sv:49:5
	output wire mem_req_rw;
	// Trace: src/VX_mem_scheduler.sv:50:5
	output wire [MEM_CHANNELS - 1:0] mem_req_mask;
	// Trace: src/VX_mem_scheduler.sv:51:5
	output wire [(MEM_CHANNELS * LINE_SIZE) - 1:0] mem_req_byteen;
	// Trace: src/VX_mem_scheduler.sv:52:5
	output wire [(MEM_CHANNELS * MEM_ADDR_WIDTH) - 1:0] mem_req_addr;
	// Trace: src/VX_mem_scheduler.sv:53:5
	output wire [(MEM_CHANNELS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] mem_req_flags;
	// Trace: src/VX_mem_scheduler.sv:54:5
	output wire [(MEM_CHANNELS * LINE_WIDTH) - 1:0] mem_req_data;
	// Trace: src/VX_mem_scheduler.sv:55:5
	output wire [MEM_TAG_WIDTH - 1:0] mem_req_tag;
	// Trace: src/VX_mem_scheduler.sv:56:5
	input wire mem_req_ready;
	// Trace: src/VX_mem_scheduler.sv:57:5
	input wire mem_rsp_valid;
	// Trace: src/VX_mem_scheduler.sv:58:5
	input wire [MEM_CHANNELS - 1:0] mem_rsp_mask;
	// Trace: src/VX_mem_scheduler.sv:59:5
	input wire [(MEM_CHANNELS * LINE_WIDTH) - 1:0] mem_rsp_data;
	// Trace: src/VX_mem_scheduler.sv:60:5
	input wire [MEM_TAG_WIDTH - 1:0] mem_rsp_tag;
	// Trace: src/VX_mem_scheduler.sv:61:5
	output wire mem_rsp_ready;
	// Trace: src/VX_mem_scheduler.sv:63:5
	localparam BATCH_SEL_WIDTH = (MEM_BATCH_BITS > 0 ? MEM_BATCH_BITS : 1);
	// Trace: src/VX_mem_scheduler.sv:64:5
	localparam STALL_TIMEOUT = 10000000;
	// Trace: src/VX_mem_scheduler.sv:65:5
	localparam TAG_ID_WIDTH = TAG_WIDTH - UUID_WIDTH;
	// Trace: src/VX_mem_scheduler.sv:66:5
	localparam REQQ_TAG_WIDTH = UUID_WIDTH + CORE_QUEUE_ADDRW;
	// Trace: src/VX_mem_scheduler.sv:67:5
	localparam MERGED_TAG_WIDTH = UUID_WIDTH + MEM_QUEUE_ADDRW;
	// Trace: src/VX_mem_scheduler.sv:68:5
	localparam CORE_CHANNELS = (COALESCE_ENABLE ? CORE_REQS : MEM_CHANNELS);
	// Trace: src/VX_mem_scheduler.sv:69:5
	localparam CORE_BATCHES = (COALESCE_ENABLE ? 1 : MEM_BATCHES);
	// Trace: src/VX_mem_scheduler.sv:70:5
	localparam CORE_BATCH_BITS = $clog2(CORE_BATCHES);
	// Trace: src/VX_mem_scheduler.sv:71:5
	wire ibuf_push;
	// Trace: src/VX_mem_scheduler.sv:72:5
	wire ibuf_pop;
	// Trace: src/VX_mem_scheduler.sv:73:5
	wire [CORE_QUEUE_ADDRW - 1:0] ibuf_waddr;
	// Trace: src/VX_mem_scheduler.sv:74:5
	wire [CORE_QUEUE_ADDRW - 1:0] ibuf_raddr;
	// Trace: src/VX_mem_scheduler.sv:75:5
	wire ibuf_full;
	// Trace: src/VX_mem_scheduler.sv:76:5
	wire ibuf_empty;
	// Trace: src/VX_mem_scheduler.sv:77:5
	wire [TAG_ID_WIDTH - 1:0] ibuf_din;
	// Trace: src/VX_mem_scheduler.sv:78:5
	wire [TAG_ID_WIDTH - 1:0] ibuf_dout;
	// Trace: src/VX_mem_scheduler.sv:79:5
	wire reqq_valid;
	// Trace: src/VX_mem_scheduler.sv:80:5
	wire [CORE_REQS - 1:0] reqq_mask;
	// Trace: src/VX_mem_scheduler.sv:81:5
	wire reqq_rw;
	// Trace: src/VX_mem_scheduler.sv:82:5
	wire [(CORE_REQS * WORD_SIZE) - 1:0] reqq_byteen;
	// Trace: src/VX_mem_scheduler.sv:83:5
	wire [(CORE_REQS * ADDR_WIDTH) - 1:0] reqq_addr;
	// Trace: src/VX_mem_scheduler.sv:84:5
	wire [(CORE_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] reqq_flags;
	// Trace: src/VX_mem_scheduler.sv:85:5
	wire [(CORE_REQS * WORD_WIDTH) - 1:0] reqq_data;
	// Trace: src/VX_mem_scheduler.sv:86:5
	wire [REQQ_TAG_WIDTH - 1:0] reqq_tag;
	// Trace: src/VX_mem_scheduler.sv:87:5
	wire reqq_ready;
	// Trace: src/VX_mem_scheduler.sv:88:5
	wire reqq_valid_s;
	// Trace: src/VX_mem_scheduler.sv:89:5
	wire [MERGED_REQS - 1:0] reqq_mask_s;
	// Trace: src/VX_mem_scheduler.sv:90:5
	wire reqq_rw_s;
	// Trace: src/VX_mem_scheduler.sv:91:5
	wire [(MERGED_REQS * LINE_SIZE) - 1:0] reqq_byteen_s;
	// Trace: src/VX_mem_scheduler.sv:92:5
	wire [(MERGED_REQS * MEM_ADDR_WIDTH) - 1:0] reqq_addr_s;
	// Trace: src/VX_mem_scheduler.sv:93:5
	wire [(MERGED_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] reqq_flags_s;
	// Trace: src/VX_mem_scheduler.sv:94:5
	wire [(MERGED_REQS * LINE_WIDTH) - 1:0] reqq_data_s;
	// Trace: src/VX_mem_scheduler.sv:95:5
	wire [MERGED_TAG_WIDTH - 1:0] reqq_tag_s;
	// Trace: src/VX_mem_scheduler.sv:96:5
	wire reqq_ready_s;
	// Trace: src/VX_mem_scheduler.sv:97:5
	wire mem_req_valid_s;
	// Trace: src/VX_mem_scheduler.sv:98:5
	wire [MEM_CHANNELS - 1:0] mem_req_mask_s;
	// Trace: src/VX_mem_scheduler.sv:99:5
	wire mem_req_rw_s;
	// Trace: src/VX_mem_scheduler.sv:100:5
	wire [(MEM_CHANNELS * LINE_SIZE) - 1:0] mem_req_byteen_s;
	// Trace: src/VX_mem_scheduler.sv:101:5
	wire [(MEM_CHANNELS * MEM_ADDR_WIDTH) - 1:0] mem_req_addr_s;
	// Trace: src/VX_mem_scheduler.sv:102:5
	wire [(MEM_CHANNELS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] mem_req_flags_s;
	// Trace: src/VX_mem_scheduler.sv:103:5
	wire [(MEM_CHANNELS * LINE_WIDTH) - 1:0] mem_req_data_s;
	// Trace: src/VX_mem_scheduler.sv:104:5
	wire [MEM_TAG_WIDTH - 1:0] mem_req_tag_s;
	// Trace: src/VX_mem_scheduler.sv:105:5
	wire mem_req_ready_s;
	// Trace: src/VX_mem_scheduler.sv:106:5
	wire mem_rsp_valid_s;
	// Trace: src/VX_mem_scheduler.sv:107:5
	wire [CORE_CHANNELS - 1:0] mem_rsp_mask_s;
	// Trace: src/VX_mem_scheduler.sv:108:5
	wire [(CORE_CHANNELS * WORD_WIDTH) - 1:0] mem_rsp_data_s;
	// Trace: src/VX_mem_scheduler.sv:109:5
	wire [MEM_TAG_WIDTH - 1:0] mem_rsp_tag_s;
	// Trace: src/VX_mem_scheduler.sv:110:5
	wire mem_rsp_ready_s;
	// Trace: src/VX_mem_scheduler.sv:111:5
	wire crsp_valid;
	// Trace: src/VX_mem_scheduler.sv:112:5
	wire [CORE_REQS - 1:0] crsp_mask;
	// Trace: src/VX_mem_scheduler.sv:113:5
	wire [(CORE_REQS * WORD_WIDTH) - 1:0] crsp_data;
	// Trace: src/VX_mem_scheduler.sv:114:5
	wire [TAG_WIDTH - 1:0] crsp_tag;
	// Trace: src/VX_mem_scheduler.sv:115:5
	wire crsp_sop;
	// Trace: src/VX_mem_scheduler.sv:116:5
	wire crsp_eop;
	// Trace: src/VX_mem_scheduler.sv:117:5
	wire crsp_ready;
	// Trace: src/VX_mem_scheduler.sv:118:5
	wire req_sent_all;
	// Trace: src/VX_mem_scheduler.sv:119:5
	wire ibuf_ready = core_req_rw || ~ibuf_full;
	// Trace: src/VX_mem_scheduler.sv:120:5
	wire reqq_valid_in = core_req_valid && ibuf_ready;
	// Trace: src/VX_mem_scheduler.sv:121:5
	wire reqq_ready_in;
	// Trace: src/VX_mem_scheduler.sv:122:5
	wire [REQQ_TAG_WIDTH - 1:0] reqq_tag_u;
	// Trace: src/VX_mem_scheduler.sv:123:5
	generate
		if (UUID_WIDTH != 0) begin : g_reqq_tag_u_uuid
			// Trace: src/VX_mem_scheduler.sv:124:9
			assign reqq_tag_u = {core_req_tag[TAG_WIDTH - 1-:UUID_WIDTH], ibuf_waddr};
		end
		else begin : g_reqq_tag_u
			// Trace: src/VX_mem_scheduler.sv:126:9
			assign reqq_tag_u = ibuf_waddr;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:128:5
	VX_elastic_buffer #(
		.DATAW((1 + (CORE_REQS * ((((1 + WORD_SIZE) + ADDR_WIDTH) + (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) + WORD_WIDTH))) + REQQ_TAG_WIDTH),
		.SIZE(CORE_QUEUE_SIZE),
		.OUT_REG(1)
	) req_queue(
		.clk(clk),
		.reset(reset),
		.valid_in(reqq_valid_in),
		.ready_in(reqq_ready_in),
		.data_in({core_req_rw, core_req_mask, core_req_byteen, core_req_addr, core_req_flags, core_req_data, reqq_tag_u}),
		.data_out({reqq_rw, reqq_mask, reqq_byteen, reqq_addr, reqq_flags, reqq_data, reqq_tag}),
		.valid_out(reqq_valid),
		.ready_out(reqq_ready)
	);
	// Trace: src/VX_mem_scheduler.sv:142:5
	assign core_req_ready = reqq_ready_in && ibuf_ready;
	// Trace: src/VX_mem_scheduler.sv:143:5
	assign req_queue_rw_notify = (reqq_valid && reqq_ready) && reqq_rw;
	// Trace: src/VX_mem_scheduler.sv:144:5
	assign req_queue_empty = !reqq_valid && ibuf_empty;
	// Trace: src/VX_mem_scheduler.sv:145:5
	wire core_req_fire = core_req_valid && core_req_ready;
	// Trace: src/VX_mem_scheduler.sv:146:5
	wire crsp_fire = crsp_valid && crsp_ready;
	// Trace: src/VX_mem_scheduler.sv:147:5
	assign ibuf_push = core_req_fire && ~core_req_rw;
	// Trace: src/VX_mem_scheduler.sv:148:5
	assign ibuf_pop = crsp_fire && crsp_eop;
	// Trace: src/VX_mem_scheduler.sv:149:5
	assign ibuf_raddr = mem_rsp_tag_s[CORE_BATCH_BITS+:CORE_QUEUE_ADDRW];
	// Trace: src/VX_mem_scheduler.sv:150:5
	assign ibuf_din = core_req_tag[TAG_ID_WIDTH - 1:0];
	// Trace: src/VX_mem_scheduler.sv:151:5
	VX_index_buffer #(
		.DATAW(TAG_ID_WIDTH),
		.SIZE(CORE_QUEUE_SIZE)
	) req_ibuf(
		.clk(clk),
		.reset(reset),
		.acquire_en(ibuf_push),
		.write_addr(ibuf_waddr),
		.write_data(ibuf_din),
		.read_data(ibuf_dout),
		.read_addr(ibuf_raddr),
		.release_en(ibuf_pop),
		.full(ibuf_full),
		.empty(ibuf_empty)
	);
	// Trace: src/VX_mem_scheduler.sv:166:5
	generate
		if (COALESCE_ENABLE) begin : g_coalescer
			// Trace: src/VX_mem_scheduler.sv:167:9
			VX_mem_coalescer #(
				.INSTANCE_ID(""),
				.NUM_REQS(CORE_REQS),
				.DATA_IN_SIZE(WORD_SIZE),
				.DATA_OUT_SIZE(LINE_SIZE),
				.ADDR_WIDTH(ADDR_WIDTH),
				.FLAGS_WIDTH(FLAGS_WIDTH),
				.TAG_WIDTH(REQQ_TAG_WIDTH),
				.UUID_WIDTH(UUID_WIDTH),
				.QUEUE_SIZE(MEM_QUEUE_SIZE)
			) coalescer(
				.clk(clk),
				.reset(reset),
				.misses(),
				.in_req_valid(reqq_valid),
				.in_req_mask(reqq_mask),
				.in_req_rw(reqq_rw),
				.in_req_byteen(reqq_byteen),
				.in_req_addr(reqq_addr),
				.in_req_flags(reqq_flags),
				.in_req_data(reqq_data),
				.in_req_tag(reqq_tag),
				.in_req_ready(reqq_ready),
				.in_rsp_valid(mem_rsp_valid_s),
				.in_rsp_mask(mem_rsp_mask_s),
				.in_rsp_data(mem_rsp_data_s),
				.in_rsp_tag(mem_rsp_tag_s),
				.in_rsp_ready(mem_rsp_ready_s),
				.out_req_valid(reqq_valid_s),
				.out_req_mask(reqq_mask_s),
				.out_req_rw(reqq_rw_s),
				.out_req_byteen(reqq_byteen_s),
				.out_req_addr(reqq_addr_s),
				.out_req_flags(reqq_flags_s),
				.out_req_data(reqq_data_s),
				.out_req_tag(reqq_tag_s),
				.out_req_ready(reqq_ready_s),
				.out_rsp_valid(mem_rsp_valid),
				.out_rsp_mask(mem_rsp_mask),
				.out_rsp_data(mem_rsp_data),
				.out_rsp_tag(mem_rsp_tag),
				.out_rsp_ready(mem_rsp_ready)
			);
		end
		else begin : g_no_coalescer
			// Trace: src/VX_mem_scheduler.sv:211:9
			assign reqq_valid_s = reqq_valid;
			// Trace: src/VX_mem_scheduler.sv:212:9
			assign reqq_mask_s = reqq_mask;
			// Trace: src/VX_mem_scheduler.sv:213:9
			assign reqq_rw_s = reqq_rw;
			// Trace: src/VX_mem_scheduler.sv:214:9
			assign reqq_byteen_s = reqq_byteen;
			// Trace: src/VX_mem_scheduler.sv:215:9
			assign reqq_addr_s = reqq_addr;
			// Trace: src/VX_mem_scheduler.sv:216:9
			assign reqq_flags_s = reqq_flags;
			// Trace: src/VX_mem_scheduler.sv:217:9
			assign reqq_data_s = reqq_data;
			// Trace: src/VX_mem_scheduler.sv:218:9
			assign reqq_tag_s = reqq_tag;
			// Trace: src/VX_mem_scheduler.sv:219:9
			assign reqq_ready = reqq_ready_s;
			// Trace: src/VX_mem_scheduler.sv:220:9
			assign mem_rsp_valid_s = mem_rsp_valid;
			// Trace: src/VX_mem_scheduler.sv:221:9
			assign mem_rsp_mask_s = mem_rsp_mask;
			// Trace: src/VX_mem_scheduler.sv:222:9
			assign mem_rsp_data_s = mem_rsp_data;
			// Trace: src/VX_mem_scheduler.sv:223:9
			assign mem_rsp_tag_s = mem_rsp_tag;
			// Trace: src/VX_mem_scheduler.sv:224:9
			assign mem_rsp_ready = mem_rsp_ready_s;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:226:5
	wire [(MEM_BATCHES * MEM_CHANNELS) - 1:0] mem_req_mask_b;
	// Trace: src/VX_mem_scheduler.sv:227:5
	wire [((MEM_BATCHES * MEM_CHANNELS) * LINE_SIZE) - 1:0] mem_req_byteen_b;
	// Trace: src/VX_mem_scheduler.sv:228:5
	wire [((MEM_BATCHES * MEM_CHANNELS) * MEM_ADDR_WIDTH) - 1:0] mem_req_addr_b;
	// Trace: src/VX_mem_scheduler.sv:229:5
	wire [((MEM_BATCHES * MEM_CHANNELS) * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] mem_req_flags_b;
	// Trace: src/VX_mem_scheduler.sv:230:5
	wire [((MEM_BATCHES * MEM_CHANNELS) * LINE_WIDTH) - 1:0] mem_req_data_b;
	// Trace: src/VX_mem_scheduler.sv:231:5
	wire [BATCH_SEL_WIDTH - 1:0] req_batch_idx;
	// Trace: src/VX_mem_scheduler.sv:232:5
	genvar _gv_i_52;
	generate
		for (_gv_i_52 = 0; _gv_i_52 < MEM_BATCHES; _gv_i_52 = _gv_i_52 + 1) begin : g_mem_req_data_b
			localparam i = _gv_i_52;
			genvar _gv_j_4;
			for (_gv_j_4 = 0; _gv_j_4 < MEM_CHANNELS; _gv_j_4 = _gv_j_4 + 1) begin : g_j
				localparam j = _gv_j_4;
				// Trace: src/VX_mem_scheduler.sv:234:13
				localparam r = (i * MEM_CHANNELS) + j;
				if (r < MERGED_REQS) begin : g_valid
					// Trace: src/VX_mem_scheduler.sv:236:17
					assign mem_req_mask_b[(i * MEM_CHANNELS) + j] = reqq_mask_s[r];
					// Trace: src/VX_mem_scheduler.sv:237:17
					assign mem_req_byteen_b[((i * MEM_CHANNELS) + j) * LINE_SIZE+:LINE_SIZE] = reqq_byteen_s[r * LINE_SIZE+:LINE_SIZE];
					// Trace: src/VX_mem_scheduler.sv:238:17
					assign mem_req_addr_b[((i * MEM_CHANNELS) + j) * MEM_ADDR_WIDTH+:MEM_ADDR_WIDTH] = reqq_addr_s[r * MEM_ADDR_WIDTH+:MEM_ADDR_WIDTH];
					// Trace: src/VX_mem_scheduler.sv:239:17
					assign mem_req_flags_b[((i * MEM_CHANNELS) + j) * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)] = reqq_flags_s[r * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)];
					// Trace: src/VX_mem_scheduler.sv:240:17
					assign mem_req_data_b[((i * MEM_CHANNELS) + j) * LINE_WIDTH+:LINE_WIDTH] = reqq_data_s[r * LINE_WIDTH+:LINE_WIDTH];
				end
				else begin : g_padding
					// Trace: src/VX_mem_scheduler.sv:242:17
					assign mem_req_mask_b[(i * MEM_CHANNELS) + j] = 0;
					// Trace: src/VX_mem_scheduler.sv:243:17
					assign mem_req_byteen_b[((i * MEM_CHANNELS) + j) * LINE_SIZE+:LINE_SIZE] = 1'sb0;
					// Trace: src/VX_mem_scheduler.sv:244:17
					assign mem_req_addr_b[((i * MEM_CHANNELS) + j) * MEM_ADDR_WIDTH+:MEM_ADDR_WIDTH] = 1'sb0;
					// Trace: src/VX_mem_scheduler.sv:245:17
					assign mem_req_flags_b[((i * MEM_CHANNELS) + j) * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)] = 1'sb0;
					// Trace: src/VX_mem_scheduler.sv:246:17
					assign mem_req_data_b[((i * MEM_CHANNELS) + j) * LINE_WIDTH+:LINE_WIDTH] = 1'sb0;
				end
			end
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:250:5
	assign mem_req_mask_s = mem_req_mask_b[req_batch_idx * MEM_CHANNELS+:MEM_CHANNELS];
	// Trace: src/VX_mem_scheduler.sv:251:5
	assign mem_req_rw_s = reqq_rw_s;
	// Trace: src/VX_mem_scheduler.sv:252:5
	assign mem_req_byteen_s = mem_req_byteen_b[LINE_SIZE * (req_batch_idx * MEM_CHANNELS)+:LINE_SIZE * MEM_CHANNELS];
	// Trace: src/VX_mem_scheduler.sv:253:5
	assign mem_req_addr_s = mem_req_addr_b[MEM_ADDR_WIDTH * (req_batch_idx * MEM_CHANNELS)+:MEM_ADDR_WIDTH * MEM_CHANNELS];
	// Trace: src/VX_mem_scheduler.sv:254:5
	assign mem_req_flags_s = mem_req_flags_b[(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1) * (req_batch_idx * MEM_CHANNELS)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1) * MEM_CHANNELS];
	// Trace: src/VX_mem_scheduler.sv:255:5
	assign mem_req_data_s = mem_req_data_b[LINE_WIDTH * (req_batch_idx * MEM_CHANNELS)+:LINE_WIDTH * MEM_CHANNELS];
	// Trace: src/VX_mem_scheduler.sv:256:5
	function automatic signed [MEM_BATCH_BITS - 1:0] sv2v_cast_F385D_signed;
		input reg signed [MEM_BATCH_BITS - 1:0] inp;
		sv2v_cast_F385D_signed = inp;
	endfunction
	generate
		if (MEM_BATCHES != 1) begin : g_batch
			// Trace: src/VX_mem_scheduler.sv:257:9
			reg [MEM_BATCH_BITS - 1:0] req_batch_idx_r;
			// Trace: src/VX_mem_scheduler.sv:258:9
			wire is_degenerate_batch = ~(|mem_req_mask_s);
			// Trace: src/VX_mem_scheduler.sv:259:9
			wire mem_req_valid_b = reqq_valid_s && ~is_degenerate_batch;
			// Trace: src/VX_mem_scheduler.sv:260:9
			wire mem_req_ready_b = mem_req_ready_s || is_degenerate_batch;
			// Trace: src/VX_mem_scheduler.sv:261:9
			always @(posedge clk)
				// Trace: src/VX_mem_scheduler.sv:262:13
				if (reset)
					// Trace: src/VX_mem_scheduler.sv:263:17
					req_batch_idx_r <= 1'sb0;
				else
					// Trace: src/VX_mem_scheduler.sv:265:17
					if (reqq_valid_s && mem_req_ready_b) begin
						begin
							// Trace: src/VX_mem_scheduler.sv:266:21
							if (req_sent_all)
								// Trace: src/VX_mem_scheduler.sv:267:25
								req_batch_idx_r <= 1'sb0;
							else
								// Trace: src/VX_mem_scheduler.sv:269:25
								req_batch_idx_r <= req_batch_idx_r + sv2v_cast_F385D_signed(1);
						end
					end
			// Trace: src/VX_mem_scheduler.sv:274:9
			wire [MEM_BATCHES - 1:0] req_batch_valids;
			// Trace: src/VX_mem_scheduler.sv:275:9
			wire [(MEM_BATCHES * MEM_BATCH_BITS) - 1:0] req_batch_idxs;
			// Trace: src/VX_mem_scheduler.sv:276:9
			wire [MEM_BATCH_BITS - 1:0] req_batch_idx_last;
			genvar _gv_i_53;
			for (_gv_i_53 = 0; _gv_i_53 < MEM_BATCHES; _gv_i_53 = _gv_i_53 + 1) begin : g_req_batch
				localparam i = _gv_i_53;
				// Trace: src/VX_mem_scheduler.sv:278:13
				assign req_batch_valids[i] = |mem_req_mask_b[i * MEM_CHANNELS+:MEM_CHANNELS];
				// Trace: src/VX_mem_scheduler.sv:279:13
				assign req_batch_idxs[i * MEM_BATCH_BITS+:MEM_BATCH_BITS] = sv2v_cast_F385D_signed(i);
			end
			// Trace: src/VX_mem_scheduler.sv:281:9
			VX_find_first #(
				.N(MEM_BATCHES),
				.DATAW(MEM_BATCH_BITS),
				.REVERSE(1)
			) find_last(
				.valid_in(req_batch_valids),
				.data_in(req_batch_idxs),
				.data_out(req_batch_idx_last),
				.valid_out()
			);
			// Trace: src/VX_mem_scheduler.sv:291:9
			assign mem_req_valid_s = mem_req_valid_b;
			// Trace: src/VX_mem_scheduler.sv:292:9
			assign req_batch_idx = req_batch_idx_r;
			// Trace: src/VX_mem_scheduler.sv:293:9
			assign req_sent_all = mem_req_ready_b && (req_batch_idx_r == req_batch_idx_last);
			// Trace: src/VX_mem_scheduler.sv:294:9
			assign mem_req_tag_s = {reqq_tag_s, req_batch_idx};
		end
		else begin : g_no_batch
			// Trace: src/VX_mem_scheduler.sv:296:9
			assign mem_req_valid_s = reqq_valid_s;
			// Trace: src/VX_mem_scheduler.sv:297:9
			assign req_batch_idx = 1'sb0;
			// Trace: src/VX_mem_scheduler.sv:298:9
			assign req_sent_all = mem_req_ready_s;
			// Trace: src/VX_mem_scheduler.sv:299:9
			assign mem_req_tag_s = reqq_tag_s;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:301:5
	assign reqq_ready_s = req_sent_all;
	// Trace: src/VX_mem_scheduler.sv:302:5
	wire [(MEM_CHANNELS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] mem_req_flags_u;
	// Trace: src/VX_mem_scheduler.sv:303:5
	VX_elastic_buffer #(
		.DATAW(((MEM_CHANNELS + 1) + (MEM_CHANNELS * (((LINE_SIZE + MEM_ADDR_WIDTH) + (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) + LINE_WIDTH))) + MEM_TAG_WIDTH),
		.SIZE(((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : 2)),
		.OUT_REG(((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : (MEM_OUT_BUF & 7) - 2))
	) mem_req_buf(
		.clk(clk),
		.reset(reset),
		.valid_in(mem_req_valid_s),
		.ready_in(mem_req_ready_s),
		.data_in({mem_req_mask_s, mem_req_rw_s, mem_req_byteen_s, mem_req_addr_s, mem_req_flags_s, mem_req_data_s, mem_req_tag_s}),
		.data_out({mem_req_mask, mem_req_rw, mem_req_byteen, mem_req_addr, mem_req_flags_u, mem_req_data, mem_req_tag}),
		.valid_out(mem_req_valid),
		.ready_out(mem_req_ready)
	);
	// Trace: src/VX_mem_scheduler.sv:317:5
	generate
		if (FLAGS_WIDTH != 0) begin : g_mem_req_flags
			// Trace: src/VX_mem_scheduler.sv:318:9
			assign mem_req_flags = mem_req_flags_u;
		end
		else begin : g_mem_req_flags_0
			// Trace: src/VX_mem_scheduler.sv:320:9
			assign mem_req_flags = 1'sb0;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:322:5
	wire [BATCH_SEL_WIDTH - 1:0] rsp_batch_idx;
	// Trace: src/VX_mem_scheduler.sv:323:5
	generate
		if (CORE_BATCHES > 1) begin : g_rsp_batch_idx
			// Trace: src/VX_mem_scheduler.sv:324:9
			assign rsp_batch_idx = mem_rsp_tag_s[CORE_BATCH_BITS - 1:0];
		end
		else begin : g_rsp_batch_idx_0
			// Trace: src/VX_mem_scheduler.sv:326:9
			assign rsp_batch_idx = 1'sb0;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:328:5
	function automatic signed [BATCH_SEL_WIDTH - 1:0] sv2v_cast_397F3_signed;
		input reg signed [BATCH_SEL_WIDTH - 1:0] inp;
		sv2v_cast_397F3_signed = inp;
	endfunction
	generate
		if (CORE_REQS == 1) begin : g_rsp_1
			// Trace: src/VX_mem_scheduler.sv:329:9
			assign crsp_valid = mem_rsp_valid_s;
			// Trace: src/VX_mem_scheduler.sv:330:9
			assign crsp_mask = mem_rsp_mask_s;
			// Trace: src/VX_mem_scheduler.sv:331:9
			assign crsp_sop = 1'b1;
			// Trace: src/VX_mem_scheduler.sv:332:9
			assign crsp_eop = 1'b1;
			// Trace: src/VX_mem_scheduler.sv:333:9
			assign crsp_data = mem_rsp_data_s;
			// Trace: src/VX_mem_scheduler.sv:334:9
			assign mem_rsp_ready_s = crsp_ready;
		end
		else begin : g_rsp_N
			// Trace: src/VX_mem_scheduler.sv:336:9
			reg [(CORE_QUEUE_SIZE * CORE_REQS) - 1:0] rsp_rem_mask;
			// Trace: src/VX_mem_scheduler.sv:337:9
			wire [CORE_REQS - 1:0] rsp_rem_mask_n;
			wire [CORE_REQS - 1:0] curr_mask;
			genvar _gv_r_1;
			for (_gv_r_1 = 0; _gv_r_1 < CORE_REQS; _gv_r_1 = _gv_r_1 + 1) begin : g_curr_mask
				localparam r = _gv_r_1;
				// Trace: src/VX_mem_scheduler.sv:339:13
				localparam i = r / CORE_CHANNELS;
				// Trace: src/VX_mem_scheduler.sv:340:13
				localparam j = r % CORE_CHANNELS;
				// Trace: src/VX_mem_scheduler.sv:341:13
				assign curr_mask[r] = (sv2v_cast_397F3_signed(i) == rsp_batch_idx) && mem_rsp_mask_s[j];
			end
			// Trace: src/VX_mem_scheduler.sv:343:9
			assign rsp_rem_mask_n = rsp_rem_mask[ibuf_raddr * CORE_REQS+:CORE_REQS] & ~curr_mask;
			// Trace: src/VX_mem_scheduler.sv:344:9
			wire mem_rsp_fire_s = mem_rsp_valid_s && mem_rsp_ready_s;
			// Trace: src/VX_mem_scheduler.sv:345:9
			always @(posedge clk) begin
				// Trace: src/VX_mem_scheduler.sv:346:13
				if (ibuf_push)
					// Trace: src/VX_mem_scheduler.sv:347:17
					rsp_rem_mask[ibuf_waddr * CORE_REQS+:CORE_REQS] <= core_req_mask;
				if (mem_rsp_fire_s)
					// Trace: src/VX_mem_scheduler.sv:350:17
					rsp_rem_mask[ibuf_raddr * CORE_REQS+:CORE_REQS] <= rsp_rem_mask_n;
			end
			// Trace: src/VX_mem_scheduler.sv:353:9
			wire rsp_complete = ~(|rsp_rem_mask_n) || (CORE_REQS == 1);
			if (RSP_PARTIAL != 0) begin : g_rsp_partial
				// Trace: src/VX_mem_scheduler.sv:355:13
				reg [CORE_QUEUE_SIZE - 1:0] rsp_sop_r;
				// Trace: src/VX_mem_scheduler.sv:356:13
				always @(posedge clk) begin
					// Trace: src/VX_mem_scheduler.sv:357:17
					if (ibuf_push)
						// Trace: src/VX_mem_scheduler.sv:358:21
						rsp_sop_r[ibuf_waddr] <= 1;
					if (mem_rsp_fire_s)
						// Trace: src/VX_mem_scheduler.sv:361:21
						rsp_sop_r[ibuf_raddr] <= 0;
				end
				// Trace: src/VX_mem_scheduler.sv:364:13
				assign crsp_valid = mem_rsp_valid_s;
				// Trace: src/VX_mem_scheduler.sv:365:13
				assign crsp_mask = curr_mask;
				// Trace: src/VX_mem_scheduler.sv:366:13
				assign crsp_sop = rsp_sop_r[ibuf_raddr];
				genvar _gv_r_2;
				for (_gv_r_2 = 0; _gv_r_2 < CORE_REQS; _gv_r_2 = _gv_r_2 + 1) begin : g_crsp_data
					localparam r = _gv_r_2;
					// Trace: src/VX_mem_scheduler.sv:368:17
					localparam j = r % CORE_CHANNELS;
					// Trace: src/VX_mem_scheduler.sv:369:17
					assign crsp_data[r * WORD_WIDTH+:WORD_WIDTH] = mem_rsp_data_s[j * WORD_WIDTH+:WORD_WIDTH];
				end
				// Trace: src/VX_mem_scheduler.sv:371:13
				assign mem_rsp_ready_s = crsp_ready;
			end
			else begin : g_rsp_full
				// Trace: src/VX_mem_scheduler.sv:373:13
				wire [((CORE_CHANNELS * CORE_BATCHES) * WORD_WIDTH) - 1:0] rsp_store_n;
				// Trace: src/VX_mem_scheduler.sv:374:13
				reg [CORE_REQS - 1:0] rsp_orig_mask [CORE_QUEUE_SIZE - 1:0];
				genvar _gv_i_54;
				for (_gv_i_54 = 0; _gv_i_54 < CORE_CHANNELS; _gv_i_54 = _gv_i_54 + 1) begin : g_rsp_store
					localparam i = _gv_i_54;
					genvar _gv_j_5;
					for (_gv_j_5 = 0; _gv_j_5 < CORE_BATCHES; _gv_j_5 = _gv_j_5 + 1) begin : g_j
						localparam j = _gv_j_5;
						// Trace: src/VX_mem_scheduler.sv:377:21
						reg [WORD_WIDTH - 1:0] rsp_store [0:CORE_QUEUE_SIZE - 1];
						// Trace: src/VX_mem_scheduler.sv:378:21
						wire rsp_wren = (mem_rsp_fire_s && (sv2v_cast_397F3_signed(j) == rsp_batch_idx)) && ((CORE_CHANNELS == 1) || mem_rsp_mask_s[i]);
						// Trace: src/VX_mem_scheduler.sv:381:21
						always @(posedge clk)
							// Trace: src/VX_mem_scheduler.sv:382:25
							if (rsp_wren)
								// Trace: src/VX_mem_scheduler.sv:383:29
								rsp_store[ibuf_raddr] <= mem_rsp_data_s[i * WORD_WIDTH+:WORD_WIDTH];
						// Trace: src/VX_mem_scheduler.sv:386:21
						assign rsp_store_n[((i * CORE_BATCHES) + j) * WORD_WIDTH+:WORD_WIDTH] = (rsp_wren ? mem_rsp_data_s[i * WORD_WIDTH+:WORD_WIDTH] : rsp_store[ibuf_raddr]);
					end
				end
				// Trace: src/VX_mem_scheduler.sv:389:13
				always @(posedge clk)
					// Trace: src/VX_mem_scheduler.sv:390:17
					if (ibuf_push)
						// Trace: src/VX_mem_scheduler.sv:391:21
						rsp_orig_mask[ibuf_waddr] <= core_req_mask;
				// Trace: src/VX_mem_scheduler.sv:394:13
				assign crsp_valid = mem_rsp_valid_s && rsp_complete;
				// Trace: src/VX_mem_scheduler.sv:395:13
				assign crsp_mask = rsp_orig_mask[ibuf_raddr];
				// Trace: src/VX_mem_scheduler.sv:396:13
				assign crsp_sop = 1'b1;
				genvar _gv_r_3;
				for (_gv_r_3 = 0; _gv_r_3 < CORE_REQS; _gv_r_3 = _gv_r_3 + 1) begin : g_crsp_data
					localparam r = _gv_r_3;
					// Trace: src/VX_mem_scheduler.sv:398:17
					localparam i = r / CORE_CHANNELS;
					// Trace: src/VX_mem_scheduler.sv:399:17
					localparam j = r % CORE_CHANNELS;
					// Trace: src/VX_mem_scheduler.sv:400:17
					assign crsp_data[r * WORD_WIDTH+:WORD_WIDTH] = rsp_store_n[((j * CORE_BATCHES) + i) * WORD_WIDTH+:WORD_WIDTH];
				end
				// Trace: src/VX_mem_scheduler.sv:402:13
				assign mem_rsp_ready_s = crsp_ready || ~rsp_complete;
			end
			// Trace: src/VX_mem_scheduler.sv:404:9
			assign crsp_eop = rsp_complete;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:406:5
	generate
		if (UUID_WIDTH != 0) begin : g_crsp_tag
			// Trace: src/VX_mem_scheduler.sv:407:9
			assign crsp_tag = {mem_rsp_tag_s[MEM_TAG_WIDTH - 1-:UUID_WIDTH], ibuf_dout};
		end
		else begin : g_crsp_tag_0
			// Trace: src/VX_mem_scheduler.sv:409:9
			assign crsp_tag = ibuf_dout;
		end
	endgenerate
	// Trace: src/VX_mem_scheduler.sv:411:5
	VX_elastic_buffer #(
		.DATAW(((CORE_REQS + 2) + (CORE_REQS * WORD_WIDTH)) + TAG_WIDTH),
		.SIZE(((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : 2)),
		.OUT_REG(((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : (CORE_OUT_BUF & 7) - 2))
	) rsp_buf(
		.clk(clk),
		.reset(reset),
		.valid_in(crsp_valid),
		.ready_in(crsp_ready),
		.data_in({crsp_mask, crsp_sop, crsp_eop, crsp_data, crsp_tag}),
		.data_out({core_rsp_mask, core_rsp_sop, core_rsp_eop, core_rsp_data, core_rsp_tag}),
		.valid_out(core_rsp_valid),
		.ready_out(core_rsp_ready)
	);
endmodule
module VX_stream_buffer (
	clk,
	reset,
	valid_in,
	ready_in,
	data_in,
	data_out,
	ready_out,
	valid_out
);
	// Trace: src/VX_stream_buffer.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_stream_buffer.sv:3:12
	parameter OUT_REG = 0;
	// Trace: src/VX_stream_buffer.sv:4:15
	parameter PASSTHRU = 0;
	// Trace: src/VX_stream_buffer.sv:6:5
	input wire clk;
	// Trace: src/VX_stream_buffer.sv:7:5
	input wire reset;
	// Trace: src/VX_stream_buffer.sv:8:5
	input wire valid_in;
	// Trace: src/VX_stream_buffer.sv:9:5
	output wire ready_in;
	// Trace: src/VX_stream_buffer.sv:10:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_stream_buffer.sv:11:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_stream_buffer.sv:12:5
	input wire ready_out;
	// Trace: src/VX_stream_buffer.sv:13:5
	output wire valid_out;
	// Trace: src/VX_stream_buffer.sv:15:5
	generate
		if (PASSTHRU != 0) begin : g_passthru
			// Trace: src/VX_stream_buffer.sv:16:9
			assign ready_in = ready_out;
			// Trace: src/VX_stream_buffer.sv:17:9
			assign valid_out = valid_in;
			// Trace: src/VX_stream_buffer.sv:18:9
			assign data_out = data_in;
		end
		else begin : g_buffer
			// Trace: src/VX_stream_buffer.sv:20:3
			reg [DATAW - 1:0] data_out_r;
			reg [DATAW - 1:0] buffer_r;
			// Trace: src/VX_stream_buffer.sv:21:3
			reg valid_out_r;
			reg valid_in_r;
			// Trace: src/VX_stream_buffer.sv:22:3
			wire fire_in = valid_in && ready_in;
			// Trace: src/VX_stream_buffer.sv:23:3
			wire flow_out = ready_out || ~valid_out;
			// Trace: src/VX_stream_buffer.sv:24:3
			always @(posedge clk)
				// Trace: src/VX_stream_buffer.sv:25:4
				if (reset)
					// Trace: src/VX_stream_buffer.sv:26:5
					valid_in_r <= 1'b1;
				else if (valid_in || flow_out)
					// Trace: src/VX_stream_buffer.sv:28:5
					valid_in_r <= flow_out;
			// Trace: src/VX_stream_buffer.sv:31:3
			always @(posedge clk)
				// Trace: src/VX_stream_buffer.sv:32:4
				if (reset)
					// Trace: src/VX_stream_buffer.sv:33:5
					valid_out_r <= 1'b0;
				else if (flow_out)
					// Trace: src/VX_stream_buffer.sv:35:5
					valid_out_r <= valid_in || ~valid_in_r;
			if (OUT_REG != 0) begin : g_out_reg
				// Trace: src/VX_stream_buffer.sv:39:4
				always @(posedge clk)
					// Trace: src/VX_stream_buffer.sv:40:5
					if (fire_in)
						// Trace: src/VX_stream_buffer.sv:41:6
						buffer_r <= data_in;
				// Trace: src/VX_stream_buffer.sv:44:4
				always @(posedge clk)
					// Trace: src/VX_stream_buffer.sv:45:5
					if (flow_out)
						// Trace: src/VX_stream_buffer.sv:46:6
						data_out_r <= (valid_in_r ? data_in : buffer_r);
				// Trace: src/VX_stream_buffer.sv:49:4
				assign data_out = data_out_r;
			end
			else begin : g_no_out_reg
				// Trace: src/VX_stream_buffer.sv:51:4
				always @(posedge clk)
					// Trace: src/VX_stream_buffer.sv:52:5
					if (fire_in)
						// Trace: src/VX_stream_buffer.sv:53:6
						data_out_r <= data_in;
				// Trace: src/VX_stream_buffer.sv:56:4
				always @(posedge clk)
					// Trace: src/VX_stream_buffer.sv:57:5
					if (fire_in)
						// Trace: src/VX_stream_buffer.sv:58:6
						buffer_r <= data_out_r;
				// Trace: src/VX_stream_buffer.sv:61:4
				assign data_out = (valid_in_r ? data_out_r : buffer_r);
			end
			// Trace: src/VX_stream_buffer.sv:63:3
			assign valid_out = valid_out_r;
			// Trace: src/VX_stream_buffer.sv:64:3
			assign ready_in = valid_in_r;
		end
	endgenerate
endmodule
// removed module with interface ports: VX_cache_bypass
// removed module with interface ports: VX_gather_unit
// removed module with interface ports: VX_ibuffer
// removed interface: VX_writeback_if
// removed module with interface ports: VX_sfu_unit
module VX_onehot_encoder (
	data_in,
	data_out,
	valid_out
);
	// Trace: src/VX_onehot_encoder.sv:2:15
	parameter N = 1;
	// Trace: src/VX_onehot_encoder.sv:3:15
	parameter REVERSE = 0;
	// Trace: src/VX_onehot_encoder.sv:4:15
	parameter MODEL = 1;
	// Trace: src/VX_onehot_encoder.sv:5:15
	parameter LN = (N > 1 ? $clog2(N) : 1);
	// Trace: src/VX_onehot_encoder.sv:7:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_onehot_encoder.sv:8:5
	output wire [LN - 1:0] data_out;
	// Trace: src/VX_onehot_encoder.sv:9:5
	output wire valid_out;
	// Trace: src/VX_onehot_encoder.sv:11:5
	function automatic signed [LN - 1:0] sv2v_cast_83428_signed;
		input reg signed [LN - 1:0] inp;
		sv2v_cast_83428_signed = inp;
	endfunction
	generate
		if (N == 1) begin : g_n1
			// Trace: src/VX_onehot_encoder.sv:12:9
			assign data_out = 0;
			// Trace: src/VX_onehot_encoder.sv:13:9
			assign valid_out = data_in;
		end
		else if (N == 2) begin : g_n2
			// Trace: src/VX_onehot_encoder.sv:15:9
			assign data_out = data_in[!REVERSE];
			// Trace: src/VX_onehot_encoder.sv:16:9
			assign valid_out = |data_in;
		end
		else if (MODEL == 1) begin : g_model1
			// Trace: src/VX_onehot_encoder.sv:18:9
			localparam M = 1 << LN;
			// Trace: src/VX_onehot_encoder.sv:19:9
			wire [M - 1:0] addr [0:LN - 1];
			// Trace: src/VX_onehot_encoder.sv:20:9
			wire [M - 1:0] v [0:LN + 0];
			// Trace: src/VX_onehot_encoder.sv:21:9
			function automatic [M - 1:0] sv2v_cast_ABEB2;
				input reg [M - 1:0] inp;
				sv2v_cast_ABEB2 = inp;
			endfunction
			assign v[0] = (REVERSE ? sv2v_cast_ABEB2(data_in) << (M - N) : sv2v_cast_ABEB2(data_in));
			genvar _gv_lvl_1;
			for (_gv_lvl_1 = 1; _gv_lvl_1 < (LN + 1); _gv_lvl_1 = _gv_lvl_1 + 1) begin : g_scan_l
				localparam lvl = _gv_lvl_1;
				// Trace: src/VX_onehot_encoder.sv:23:13
				localparam SN = 1 << (LN - lvl);
				// Trace: src/VX_onehot_encoder.sv:24:13
				localparam SI = M / SN;
				genvar _gv_s_1;
				for (_gv_s_1 = 0; _gv_s_1 < SN; _gv_s_1 = _gv_s_1 + 1) begin : g_scan_s
					localparam s = _gv_s_1;
					// Trace: src/VX_onehot_encoder.sv:26:17
					wire [1:0] vs = {v[lvl - 1][(s * SI) + (SI >> 1)], v[lvl - 1][s * SI]};
					// Trace: src/VX_onehot_encoder.sv:27:17
					assign v[lvl][s * SI] = |vs;
					if (lvl == 1) begin : g_lvl_1
						// Trace: src/VX_onehot_encoder.sv:29:21
						assign addr[lvl - 1][s * SI+:lvl] = vs[!REVERSE];
					end
					else begin : g_lvl_n
						// Trace: src/VX_onehot_encoder.sv:31:21
						assign addr[lvl - 1][s * SI+:lvl] = {vs[!REVERSE], addr[lvl - 2][s * SI+:lvl - 1] | addr[lvl - 2][(s * SI) + (SI >> 1)+:lvl - 1]};
					end
				end
			end
			// Trace: src/VX_onehot_encoder.sv:38:9
			assign data_out = addr[LN - 1][LN - 1:0];
			// Trace: src/VX_onehot_encoder.sv:39:9
			assign valid_out = v[LN][0];
		end
		else if ((MODEL == 2) && (REVERSE == 0)) begin : g_model2
			genvar _gv_j_6;
			for (_gv_j_6 = 0; _gv_j_6 < LN; _gv_j_6 = _gv_j_6 + 1) begin : g_data_out
				localparam j = _gv_j_6;
				// Trace: src/VX_onehot_encoder.sv:42:13
				wire [N - 1:0] mask;
				genvar _gv_i_66;
				for (_gv_i_66 = 0; _gv_i_66 < N; _gv_i_66 = _gv_i_66 + 1) begin : g_mask
					localparam i = _gv_i_66;
					// Trace: src/VX_onehot_encoder.sv:44:17
					assign mask[i] = i[j];
				end
				// Trace: src/VX_onehot_encoder.sv:46:13
				assign data_out[j] = |(mask & data_in);
			end
			// Trace: src/VX_onehot_encoder.sv:48:9
			assign valid_out = |data_in;
		end
		else begin : g_model0
			// Trace: src/VX_onehot_encoder.sv:50:9
			reg [LN - 1:0] index_w;
			if (REVERSE != 0) begin : g_msb
				// Trace: src/VX_onehot_encoder.sv:52:13
				always @(*) begin
					// Trace: src/VX_onehot_encoder.sv:53:17
					index_w = 1'sbx;
					// Trace: src/VX_onehot_encoder.sv:54:17
					begin : sv2v_autoblock_1
						// Trace: src/VX_onehot_encoder.sv:54:22
						integer i;
						// Trace: src/VX_onehot_encoder.sv:54:22
						for (i = N - 1; i >= 0; i = i - 1)
							begin
								// Trace: src/VX_onehot_encoder.sv:55:21
								if (data_in[i])
									// Trace: src/VX_onehot_encoder.sv:56:25
									index_w = sv2v_cast_83428_signed((N - 1) - i);
							end
					end
				end
			end
			else begin : g_lsb
				// Trace: src/VX_onehot_encoder.sv:61:13
				always @(*) begin
					// Trace: src/VX_onehot_encoder.sv:62:17
					index_w = 1'sbx;
					// Trace: src/VX_onehot_encoder.sv:63:17
					begin : sv2v_autoblock_2
						// Trace: src/VX_onehot_encoder.sv:63:22
						integer i;
						// Trace: src/VX_onehot_encoder.sv:63:22
						for (i = 0; i < N; i = i + 1)
							begin
								// Trace: src/VX_onehot_encoder.sv:64:21
								if (data_in[i])
									// Trace: src/VX_onehot_encoder.sv:65:25
									index_w = sv2v_cast_83428_signed(i);
							end
					end
				end
			end
			// Trace: src/VX_onehot_encoder.sv:70:9
			assign data_out = index_w;
			// Trace: src/VX_onehot_encoder.sv:71:9
			assign valid_out = |data_in;
		end
	endgenerate
endmodule
module VX_cache_mshr (
	clk,
	reset,
	deq_req_uuid,
	alc_req_uuid,
	fin_req_uuid,
	fill_valid,
	fill_id,
	fill_addr,
	dequeue_valid,
	dequeue_addr,
	dequeue_rw,
	dequeue_data,
	dequeue_id,
	dequeue_ready,
	allocate_valid,
	allocate_addr,
	allocate_rw,
	allocate_data,
	allocate_id,
	allocate_pending,
	allocate_previd,
	allocate_ready,
	finalize_valid,
	finalize_is_release,
	finalize_is_pending,
	finalize_previd,
	finalize_id
);
	// removed import VX_gpu_pkg::*;
	// Trace: src/VX_cache_mshr.sv:2:15
	parameter INSTANCE_ID = "";
	// Trace: src/VX_cache_mshr.sv:3:15
	parameter BANK_ID = 0;
	// Trace: src/VX_cache_mshr.sv:4:15
	parameter LINE_SIZE = 16;
	// Trace: src/VX_cache_mshr.sv:5:15
	parameter NUM_BANKS = 1;
	// Trace: src/VX_cache_mshr.sv:6:15
	parameter MSHR_SIZE = 4;
	// Trace: src/VX_cache_mshr.sv:7:15
	parameter DATA_WIDTH = 1;
	// Trace: src/VX_cache_mshr.sv:8:15
	parameter WRITEBACK = 0;
	// Trace: src/VX_cache_mshr.sv:9:15
	parameter MSHR_ADDR_WIDTH = (MSHR_SIZE > 1 ? $clog2(MSHR_SIZE) : 1);
	// Trace: src/VX_cache_mshr.sv:11:5
	input wire clk;
	// Trace: src/VX_cache_mshr.sv:12:5
	input wire reset;
	// Trace: src/VX_cache_mshr.sv:13:5
	localparam VX_gpu_pkg_UUID_WIDTH = 1;
	input wire [0:0] deq_req_uuid;
	// Trace: src/VX_cache_mshr.sv:14:5
	input wire [0:0] alc_req_uuid;
	// Trace: src/VX_cache_mshr.sv:15:5
	input wire [0:0] fin_req_uuid;
	// Trace: src/VX_cache_mshr.sv:16:5
	input wire fill_valid;
	// Trace: src/VX_cache_mshr.sv:17:5
	input wire [MSHR_ADDR_WIDTH - 1:0] fill_id;
	// Trace: src/VX_cache_mshr.sv:18:5
	output wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] fill_addr;
	// Trace: src/VX_cache_mshr.sv:19:5
	output wire dequeue_valid;
	// Trace: src/VX_cache_mshr.sv:20:5
	output wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] dequeue_addr;
	// Trace: src/VX_cache_mshr.sv:21:5
	output wire dequeue_rw;
	// Trace: src/VX_cache_mshr.sv:22:5
	output wire [DATA_WIDTH - 1:0] dequeue_data;
	// Trace: src/VX_cache_mshr.sv:23:5
	output wire [MSHR_ADDR_WIDTH - 1:0] dequeue_id;
	// Trace: src/VX_cache_mshr.sv:24:5
	input wire dequeue_ready;
	// Trace: src/VX_cache_mshr.sv:25:5
	input wire allocate_valid;
	// Trace: src/VX_cache_mshr.sv:26:5
	input wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] allocate_addr;
	// Trace: src/VX_cache_mshr.sv:27:5
	input wire allocate_rw;
	// Trace: src/VX_cache_mshr.sv:28:5
	input wire [DATA_WIDTH - 1:0] allocate_data;
	// Trace: src/VX_cache_mshr.sv:29:5
	output wire [MSHR_ADDR_WIDTH - 1:0] allocate_id;
	// Trace: src/VX_cache_mshr.sv:30:5
	output wire allocate_pending;
	// Trace: src/VX_cache_mshr.sv:31:5
	output wire [MSHR_ADDR_WIDTH - 1:0] allocate_previd;
	// Trace: src/VX_cache_mshr.sv:32:5
	output wire allocate_ready;
	// Trace: src/VX_cache_mshr.sv:33:5
	input wire finalize_valid;
	// Trace: src/VX_cache_mshr.sv:34:5
	input wire finalize_is_release;
	// Trace: src/VX_cache_mshr.sv:35:5
	input wire finalize_is_pending;
	// Trace: src/VX_cache_mshr.sv:36:5
	input wire [MSHR_ADDR_WIDTH - 1:0] finalize_previd;
	// Trace: src/VX_cache_mshr.sv:37:5
	input wire [MSHR_ADDR_WIDTH - 1:0] finalize_id;
	// Trace: src/VX_cache_mshr.sv:39:5
	reg [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] addr_table [0:MSHR_SIZE - 1];
	// Trace: src/VX_cache_mshr.sv:40:5
	reg [MSHR_ADDR_WIDTH - 1:0] next_index [0:MSHR_SIZE - 1];
	// Trace: src/VX_cache_mshr.sv:41:5
	reg [MSHR_SIZE - 1:0] valid_table;
	reg [MSHR_SIZE - 1:0] valid_table_n;
	// Trace: src/VX_cache_mshr.sv:42:5
	reg [MSHR_SIZE - 1:0] next_table;
	reg [MSHR_SIZE - 1:0] next_table_x;
	reg [MSHR_SIZE - 1:0] next_table_n;
	// Trace: src/VX_cache_mshr.sv:43:5
	reg [MSHR_SIZE - 1:0] write_table;
	// Trace: src/VX_cache_mshr.sv:44:5
	reg allocate_rdy;
	reg allocate_rdy_n;
	// Trace: src/VX_cache_mshr.sv:45:5
	reg [MSHR_ADDR_WIDTH - 1:0] allocate_id_r;
	reg [MSHR_ADDR_WIDTH - 1:0] allocate_id_n;
	// Trace: src/VX_cache_mshr.sv:46:5
	reg dequeue_val;
	reg dequeue_val_n;
	// Trace: src/VX_cache_mshr.sv:47:5
	reg [MSHR_ADDR_WIDTH - 1:0] dequeue_id_r;
	reg [MSHR_ADDR_WIDTH - 1:0] dequeue_id_n;
	// Trace: src/VX_cache_mshr.sv:48:5
	wire [MSHR_ADDR_WIDTH - 1:0] prev_idx;
	// Trace: src/VX_cache_mshr.sv:49:5
	wire allocate_fire = allocate_valid && allocate_ready;
	// Trace: src/VX_cache_mshr.sv:50:5
	wire dequeue_fire = dequeue_valid && dequeue_ready;
	// Trace: src/VX_cache_mshr.sv:51:5
	wire [MSHR_SIZE - 1:0] addr_matches;
	// Trace: src/VX_cache_mshr.sv:52:5
	genvar _gv_i_67;
	generate
		for (_gv_i_67 = 0; _gv_i_67 < MSHR_SIZE; _gv_i_67 = _gv_i_67 + 1) begin : g_addr_matches
			localparam i = _gv_i_67;
			// Trace: src/VX_cache_mshr.sv:53:9
			assign addr_matches[i] = valid_table[i] && (addr_table[i] == allocate_addr);
		end
	endgenerate
	// Trace: src/VX_cache_mshr.sv:55:5
	// rewrote reg-to-output bindings
	wire [MSHR_ADDR_WIDTH:1] sv2v_tmp_allocate_sel_index_out;
	always @(*) allocate_id_n = sv2v_tmp_allocate_sel_index_out;
	wire [1:1] sv2v_tmp_allocate_sel_valid_out;
	always @(*) allocate_rdy_n = sv2v_tmp_allocate_sel_valid_out;
	VX_priority_encoder #(.N(MSHR_SIZE)) allocate_sel(
		.data_in(~valid_table_n),
		.index_out(sv2v_tmp_allocate_sel_index_out),
		.valid_out(sv2v_tmp_allocate_sel_valid_out),
		.onehot_out()
	);
	// Trace: src/VX_cache_mshr.sv:63:5
	VX_priority_encoder #(.N(MSHR_SIZE)) prev_sel(
		.data_in(addr_matches & ~next_table_x),
		.index_out(prev_idx),
		.valid_out(),
		.onehot_out()
	);
	// Trace: src/VX_cache_mshr.sv:71:5
	always @(*) begin
		// Trace: src/VX_cache_mshr.sv:72:9
		valid_table_n = valid_table;
		// Trace: src/VX_cache_mshr.sv:73:9
		next_table_x = next_table;
		// Trace: src/VX_cache_mshr.sv:74:9
		dequeue_val_n = dequeue_val;
		// Trace: src/VX_cache_mshr.sv:75:9
		dequeue_id_n = dequeue_id;
		// Trace: src/VX_cache_mshr.sv:76:9
		if (fill_valid) begin
			// Trace: src/VX_cache_mshr.sv:77:13
			dequeue_val_n = 1;
			// Trace: src/VX_cache_mshr.sv:78:13
			dequeue_id_n = fill_id;
		end
		if (dequeue_fire) begin
			// Trace: src/VX_cache_mshr.sv:81:13
			valid_table_n[dequeue_id] = 0;
			// Trace: src/VX_cache_mshr.sv:82:13
			if (next_table[dequeue_id])
				// Trace: src/VX_cache_mshr.sv:83:17
				dequeue_id_n = next_index[dequeue_id];
			else if ((finalize_valid && finalize_is_pending) && (finalize_previd == dequeue_id))
				// Trace: src/VX_cache_mshr.sv:85:17
				dequeue_id_n = finalize_id;
			else
				// Trace: src/VX_cache_mshr.sv:87:17
				dequeue_val_n = 0;
		end
		if (finalize_valid) begin
			// Trace: src/VX_cache_mshr.sv:91:13
			if (finalize_is_release)
				// Trace: src/VX_cache_mshr.sv:92:17
				valid_table_n[finalize_id] = 0;
			if (finalize_is_pending)
				// Trace: src/VX_cache_mshr.sv:95:17
				next_table_x[finalize_previd] = 1;
		end
		// Trace: src/VX_cache_mshr.sv:98:9
		next_table_n = next_table_x;
		if (allocate_fire) begin
			// Trace: src/VX_cache_mshr.sv:100:13
			valid_table_n[allocate_id] = 1;
			// Trace: src/VX_cache_mshr.sv:101:13
			next_table_n[allocate_id] = 0;
		end
	end
	// Trace: src/VX_cache_mshr.sv:104:5
	always @(posedge clk) begin
		// Trace: src/VX_cache_mshr.sv:105:9
		if (reset) begin
			// Trace: src/VX_cache_mshr.sv:106:13
			valid_table <= 1'sb0;
			// Trace: src/VX_cache_mshr.sv:107:13
			allocate_rdy <= 0;
			// Trace: src/VX_cache_mshr.sv:108:13
			dequeue_val <= 0;
		end
		else begin
			// Trace: src/VX_cache_mshr.sv:110:13
			valid_table <= valid_table_n;
			// Trace: src/VX_cache_mshr.sv:111:13
			allocate_rdy <= allocate_rdy_n;
			// Trace: src/VX_cache_mshr.sv:112:13
			dequeue_val <= dequeue_val_n;
		end
		if (allocate_fire) begin
			// Trace: src/VX_cache_mshr.sv:115:13
			addr_table[allocate_id] <= allocate_addr;
			// Trace: src/VX_cache_mshr.sv:116:13
			write_table[allocate_id] <= allocate_rw;
		end
		if (finalize_valid && finalize_is_pending)
			// Trace: src/VX_cache_mshr.sv:119:13
			next_index[finalize_previd] <= finalize_id;
		// Trace: src/VX_cache_mshr.sv:121:9
		dequeue_id_r <= dequeue_id_n;
		// Trace: src/VX_cache_mshr.sv:122:9
		allocate_id_r <= allocate_id_n;
		// Trace: src/VX_cache_mshr.sv:123:9
		next_table <= next_table_n;
	end
	// Trace: src/VX_cache_mshr.sv:125:5
	VX_dp_ram #(
		.DATAW(DATA_WIDTH),
		.SIZE(MSHR_SIZE),
		.RDW_MODE("R"),
		.RADDR_REG(1)
	) mshr_store(
		.clk(clk),
		.reset(reset),
		.read(1'b1),
		.write(allocate_valid),
		.wren(1'b1),
		.waddr(allocate_id_r),
		.wdata(allocate_data),
		.raddr(dequeue_id_r),
		.rdata(dequeue_data)
	);
	// Trace: src/VX_cache_mshr.sv:141:5
	assign fill_addr = addr_table[fill_id];
	// Trace: src/VX_cache_mshr.sv:142:5
	assign allocate_ready = allocate_rdy;
	// Trace: src/VX_cache_mshr.sv:143:5
	assign allocate_id = allocate_id_r;
	// Trace: src/VX_cache_mshr.sv:144:5
	assign allocate_previd = prev_idx;
	// Trace: src/VX_cache_mshr.sv:145:5
	generate
		if (WRITEBACK) begin : g_pending_wb
			// Trace: src/VX_cache_mshr.sv:146:9
			assign allocate_pending = |addr_matches;
		end
		else begin : g_pending_wt
			// Trace: src/VX_cache_mshr.sv:148:9
			assign allocate_pending = |(addr_matches & ~write_table);
		end
	endgenerate
	// Trace: src/VX_cache_mshr.sv:150:5
	assign dequeue_valid = dequeue_val;
	// Trace: src/VX_cache_mshr.sv:151:5
	assign dequeue_addr = addr_table[dequeue_id_r];
	// Trace: src/VX_cache_mshr.sv:152:5
	assign dequeue_rw = write_table[dequeue_id_r];
	// Trace: src/VX_cache_mshr.sv:153:5
	assign dequeue_id = dequeue_id_r;
endmodule
module VX_mem_coalescer (
	clk,
	reset,
	misses,
	in_req_valid,
	in_req_rw,
	in_req_mask,
	in_req_byteen,
	in_req_addr,
	in_req_flags,
	in_req_data,
	in_req_tag,
	in_req_ready,
	in_rsp_valid,
	in_rsp_mask,
	in_rsp_data,
	in_rsp_tag,
	in_rsp_ready,
	out_req_valid,
	out_req_rw,
	out_req_mask,
	out_req_byteen,
	out_req_addr,
	out_req_flags,
	out_req_data,
	out_req_tag,
	out_req_ready,
	out_rsp_valid,
	out_rsp_mask,
	out_rsp_data,
	out_rsp_tag,
	out_rsp_ready
);
	// Trace: src/VX_mem_coalescer.sv:2:15
	parameter INSTANCE_ID = "";
	// Trace: src/VX_mem_coalescer.sv:3:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_mem_coalescer.sv:4:15
	parameter ADDR_WIDTH = 32;
	// Trace: src/VX_mem_coalescer.sv:5:15
	parameter FLAGS_WIDTH = 0;
	// Trace: src/VX_mem_coalescer.sv:6:15
	parameter DATA_IN_SIZE = 4;
	// Trace: src/VX_mem_coalescer.sv:7:15
	parameter DATA_OUT_SIZE = 64;
	// Trace: src/VX_mem_coalescer.sv:8:15
	parameter TAG_WIDTH = 8;
	// Trace: src/VX_mem_coalescer.sv:9:15
	parameter UUID_WIDTH = 0;
	// Trace: src/VX_mem_coalescer.sv:10:15
	parameter QUEUE_SIZE = 8;
	// Trace: src/VX_mem_coalescer.sv:11:15
	parameter PERF_CTR_BITS = $clog2(NUM_REQS + 1);
	// Trace: src/VX_mem_coalescer.sv:12:15
	parameter DATA_IN_WIDTH = DATA_IN_SIZE * 8;
	// Trace: src/VX_mem_coalescer.sv:13:15
	parameter DATA_OUT_WIDTH = DATA_OUT_SIZE * 8;
	// Trace: src/VX_mem_coalescer.sv:14:15
	parameter DATA_RATIO = DATA_OUT_SIZE / DATA_IN_SIZE;
	// Trace: src/VX_mem_coalescer.sv:15:15
	parameter DATA_RATIO_W = (DATA_RATIO > 1 ? $clog2(DATA_RATIO) : 1);
	// Trace: src/VX_mem_coalescer.sv:16:15
	parameter OUT_REQS = NUM_REQS / DATA_RATIO;
	// Trace: src/VX_mem_coalescer.sv:17:15
	parameter OUT_ADDR_WIDTH = ADDR_WIDTH - DATA_RATIO_W;
	// Trace: src/VX_mem_coalescer.sv:18:15
	parameter QUEUE_ADDRW = $clog2(QUEUE_SIZE);
	// Trace: src/VX_mem_coalescer.sv:19:15
	parameter OUT_TAG_WIDTH = UUID_WIDTH + QUEUE_ADDRW;
	// Trace: src/VX_mem_coalescer.sv:21:5
	input wire clk;
	// Trace: src/VX_mem_coalescer.sv:22:5
	input wire reset;
	// Trace: src/VX_mem_coalescer.sv:23:5
	output wire [PERF_CTR_BITS - 1:0] misses;
	// Trace: src/VX_mem_coalescer.sv:24:5
	input wire in_req_valid;
	// Trace: src/VX_mem_coalescer.sv:25:5
	input wire in_req_rw;
	// Trace: src/VX_mem_coalescer.sv:26:5
	input wire [NUM_REQS - 1:0] in_req_mask;
	// Trace: src/VX_mem_coalescer.sv:27:5
	input wire [(NUM_REQS * DATA_IN_SIZE) - 1:0] in_req_byteen;
	// Trace: src/VX_mem_coalescer.sv:28:5
	input wire [(NUM_REQS * ADDR_WIDTH) - 1:0] in_req_addr;
	// Trace: src/VX_mem_coalescer.sv:29:5
	input wire [(NUM_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] in_req_flags;
	// Trace: src/VX_mem_coalescer.sv:30:5
	input wire [(NUM_REQS * DATA_IN_WIDTH) - 1:0] in_req_data;
	// Trace: src/VX_mem_coalescer.sv:31:5
	input wire [TAG_WIDTH - 1:0] in_req_tag;
	// Trace: src/VX_mem_coalescer.sv:32:5
	output wire in_req_ready;
	// Trace: src/VX_mem_coalescer.sv:33:5
	output wire in_rsp_valid;
	// Trace: src/VX_mem_coalescer.sv:34:5
	output wire [NUM_REQS - 1:0] in_rsp_mask;
	// Trace: src/VX_mem_coalescer.sv:35:5
	output wire [(NUM_REQS * DATA_IN_WIDTH) - 1:0] in_rsp_data;
	// Trace: src/VX_mem_coalescer.sv:36:5
	output wire [TAG_WIDTH - 1:0] in_rsp_tag;
	// Trace: src/VX_mem_coalescer.sv:37:5
	input wire in_rsp_ready;
	// Trace: src/VX_mem_coalescer.sv:38:5
	output wire out_req_valid;
	// Trace: src/VX_mem_coalescer.sv:39:5
	output wire out_req_rw;
	// Trace: src/VX_mem_coalescer.sv:40:5
	output wire [OUT_REQS - 1:0] out_req_mask;
	// Trace: src/VX_mem_coalescer.sv:41:5
	output wire [(OUT_REQS * DATA_OUT_SIZE) - 1:0] out_req_byteen;
	// Trace: src/VX_mem_coalescer.sv:42:5
	output wire [(OUT_REQS * OUT_ADDR_WIDTH) - 1:0] out_req_addr;
	// Trace: src/VX_mem_coalescer.sv:43:5
	output wire [(OUT_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] out_req_flags;
	// Trace: src/VX_mem_coalescer.sv:44:5
	output wire [(OUT_REQS * DATA_OUT_WIDTH) - 1:0] out_req_data;
	// Trace: src/VX_mem_coalescer.sv:45:5
	output wire [OUT_TAG_WIDTH - 1:0] out_req_tag;
	// Trace: src/VX_mem_coalescer.sv:46:5
	input wire out_req_ready;
	// Trace: src/VX_mem_coalescer.sv:47:5
	input wire out_rsp_valid;
	// Trace: src/VX_mem_coalescer.sv:48:5
	input wire [OUT_REQS - 1:0] out_rsp_mask;
	// Trace: src/VX_mem_coalescer.sv:49:5
	input wire [(OUT_REQS * DATA_OUT_WIDTH) - 1:0] out_rsp_data;
	// Trace: src/VX_mem_coalescer.sv:50:5
	input wire [OUT_TAG_WIDTH - 1:0] out_rsp_tag;
	// Trace: src/VX_mem_coalescer.sv:51:5
	output wire out_rsp_ready;
	// Trace: src/VX_mem_coalescer.sv:53:5
	localparam TAG_ID_WIDTH = TAG_WIDTH - UUID_WIDTH;
	// Trace: src/VX_mem_coalescer.sv:54:5
	localparam IBUF_DATA_WIDTH = (TAG_ID_WIDTH + NUM_REQS) + (NUM_REQS * DATA_RATIO_W);
	// Trace: src/VX_mem_coalescer.sv:55:5
	localparam STATE_WAIT = 0;
	// Trace: src/VX_mem_coalescer.sv:56:5
	localparam STATE_SEND = 1;
	// Trace: src/VX_mem_coalescer.sv:57:5
	wire state_r;
	reg state_n;
	// Trace: src/VX_mem_coalescer.sv:58:5
	wire out_req_valid_r;
	reg out_req_valid_n;
	// Trace: src/VX_mem_coalescer.sv:59:5
	wire out_req_rw_r;
	reg out_req_rw_n;
	// Trace: src/VX_mem_coalescer.sv:60:5
	wire [OUT_REQS - 1:0] out_req_mask_r;
	reg [OUT_REQS - 1:0] out_req_mask_n;
	// Trace: src/VX_mem_coalescer.sv:61:5
	wire [(OUT_REQS * OUT_ADDR_WIDTH) - 1:0] out_req_addr_r;
	reg [(OUT_REQS * OUT_ADDR_WIDTH) - 1:0] out_req_addr_n;
	// Trace: src/VX_mem_coalescer.sv:62:5
	wire [(OUT_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] out_req_flags_r;
	reg [(OUT_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] out_req_flags_n;
	// Trace: src/VX_mem_coalescer.sv:63:5
	wire [((OUT_REQS * DATA_RATIO) * DATA_IN_SIZE) - 1:0] out_req_byteen_r;
	reg [((OUT_REQS * DATA_RATIO) * DATA_IN_SIZE) - 1:0] out_req_byteen_n;
	// Trace: src/VX_mem_coalescer.sv:64:5
	wire [((OUT_REQS * DATA_RATIO) * DATA_IN_WIDTH) - 1:0] out_req_data_r;
	reg [((OUT_REQS * DATA_RATIO) * DATA_IN_WIDTH) - 1:0] out_req_data_n;
	// Trace: src/VX_mem_coalescer.sv:65:5
	wire [OUT_TAG_WIDTH - 1:0] out_req_tag_r;
	reg [OUT_TAG_WIDTH - 1:0] out_req_tag_n;
	// Trace: src/VX_mem_coalescer.sv:66:5
	reg in_req_ready_n;
	// Trace: src/VX_mem_coalescer.sv:67:5
	wire ibuf_push;
	// Trace: src/VX_mem_coalescer.sv:68:5
	wire ibuf_pop;
	// Trace: src/VX_mem_coalescer.sv:69:5
	wire [QUEUE_ADDRW - 1:0] ibuf_waddr;
	// Trace: src/VX_mem_coalescer.sv:70:5
	wire [QUEUE_ADDRW - 1:0] ibuf_raddr;
	// Trace: src/VX_mem_coalescer.sv:71:5
	wire ibuf_full;
	// Trace: src/VX_mem_coalescer.sv:72:5
	wire ibuf_empty;
	// Trace: src/VX_mem_coalescer.sv:73:5
	wire [IBUF_DATA_WIDTH - 1:0] ibuf_din;
	// Trace: src/VX_mem_coalescer.sv:74:5
	wire [IBUF_DATA_WIDTH - 1:0] ibuf_dout;
	// Trace: src/VX_mem_coalescer.sv:75:5
	wire [OUT_REQS - 1:0] batch_valid_r;
	wire [OUT_REQS - 1:0] batch_valid_n;
	// Trace: src/VX_mem_coalescer.sv:76:5
	wire [(OUT_REQS * OUT_ADDR_WIDTH) - 1:0] seed_addr_r;
	wire [(OUT_REQS * OUT_ADDR_WIDTH) - 1:0] seed_addr_n;
	// Trace: src/VX_mem_coalescer.sv:77:5
	wire [(OUT_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] seed_flags_r;
	wire [(OUT_REQS * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] seed_flags_n;
	// Trace: src/VX_mem_coalescer.sv:78:5
	wire [NUM_REQS - 1:0] addr_matches_r;
	wire [NUM_REQS - 1:0] addr_matches_n;
	// Trace: src/VX_mem_coalescer.sv:79:5
	wire [NUM_REQS - 1:0] req_rem_mask_r;
	reg [NUM_REQS - 1:0] req_rem_mask_n;
	// Trace: src/VX_mem_coalescer.sv:80:5
	wire [(NUM_REQS * DATA_RATIO_W) - 1:0] in_addr_offset;
	// Trace: src/VX_mem_coalescer.sv:81:5
	genvar _gv_i_68;
	generate
		for (_gv_i_68 = 0; _gv_i_68 < NUM_REQS; _gv_i_68 = _gv_i_68 + 1) begin : g_in_addr_offset
			localparam i = _gv_i_68;
			// Trace: src/VX_mem_coalescer.sv:82:9
			assign in_addr_offset[i * DATA_RATIO_W+:DATA_RATIO_W] = in_req_addr[(i * ADDR_WIDTH) + (DATA_RATIO_W - 1)-:DATA_RATIO_W];
		end
	endgenerate
	// Trace: src/VX_mem_coalescer.sv:84:5
	genvar _gv_i_69;
	generate
		for (_gv_i_69 = 0; _gv_i_69 < OUT_REQS; _gv_i_69 = _gv_i_69 + 1) begin : g_seed_gen
			localparam i = _gv_i_69;
			// Trace: src/VX_mem_coalescer.sv:85:9
			wire [DATA_RATIO - 1:0] batch_mask;
			// Trace: src/VX_mem_coalescer.sv:86:9
			wire [DATA_RATIO_W - 1:0] batch_idx;
			// Trace: src/VX_mem_coalescer.sv:87:9
			assign batch_mask = in_req_mask[i * DATA_RATIO+:DATA_RATIO] & req_rem_mask_r[i * DATA_RATIO+:DATA_RATIO];
			// Trace: src/VX_mem_coalescer.sv:88:9
			VX_priority_encoder #(.N(DATA_RATIO)) batch_sel(
				.data_in(batch_mask),
				.index_out(batch_idx),
				.valid_out(batch_valid_n[i]),
				.onehot_out()
			);
			// Trace: src/VX_mem_coalescer.sv:96:9
			wire [(DATA_RATIO * OUT_ADDR_WIDTH) - 1:0] addr_base;
			genvar _gv_j_7;
			for (_gv_j_7 = 0; _gv_j_7 < DATA_RATIO; _gv_j_7 = _gv_j_7 + 1) begin : g_addr_base
				localparam j = _gv_j_7;
				// Trace: src/VX_mem_coalescer.sv:98:13
				assign addr_base[j * OUT_ADDR_WIDTH+:OUT_ADDR_WIDTH] = in_req_addr[(((DATA_RATIO * i) + j) * ADDR_WIDTH) + ((ADDR_WIDTH - 1) >= DATA_RATIO_W ? ADDR_WIDTH - 1 : ((ADDR_WIDTH - 1) + ((ADDR_WIDTH - 1) >= DATA_RATIO_W ? ((ADDR_WIDTH - 1) - DATA_RATIO_W) + 1 : (DATA_RATIO_W - (ADDR_WIDTH - 1)) + 1)) - 1)-:((ADDR_WIDTH - 1) >= DATA_RATIO_W ? ((ADDR_WIDTH - 1) - DATA_RATIO_W) + 1 : (DATA_RATIO_W - (ADDR_WIDTH - 1)) + 1)];
			end
			// Trace: src/VX_mem_coalescer.sv:100:9
			wire [(DATA_RATIO * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) - 1:0] req_flags;
			genvar _gv_j_8;
			for (_gv_j_8 = 0; _gv_j_8 < DATA_RATIO; _gv_j_8 = _gv_j_8 + 1) begin : g_req_flags
				localparam j = _gv_j_8;
				// Trace: src/VX_mem_coalescer.sv:102:13
				assign req_flags[j * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)] = in_req_flags[((DATA_RATIO * i) + j) * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)];
			end
			// Trace: src/VX_mem_coalescer.sv:104:9
			assign seed_addr_n[i * OUT_ADDR_WIDTH+:OUT_ADDR_WIDTH] = addr_base[batch_idx * OUT_ADDR_WIDTH+:OUT_ADDR_WIDTH];
			// Trace: src/VX_mem_coalescer.sv:105:9
			assign seed_flags_n[i * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)] = req_flags[batch_idx * (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)+:(FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)];
			genvar _gv_j_9;
			for (_gv_j_9 = 0; _gv_j_9 < DATA_RATIO; _gv_j_9 = _gv_j_9 + 1) begin : g_addr_matches_n
				localparam j = _gv_j_9;
				// Trace: src/VX_mem_coalescer.sv:107:13
				assign addr_matches_n[(i * DATA_RATIO) + j] = addr_base[j * OUT_ADDR_WIDTH+:OUT_ADDR_WIDTH] == seed_addr_n[i * OUT_ADDR_WIDTH+:OUT_ADDR_WIDTH];
			end
		end
	endgenerate
	// Trace: src/VX_mem_coalescer.sv:110:5
	wire [NUM_REQS - 1:0] current_pmask = in_req_mask & addr_matches_r;
	// Trace: src/VX_mem_coalescer.sv:111:5
	wire [((OUT_REQS * DATA_RATIO) * DATA_IN_SIZE) - 1:0] req_byteen_merged;
	// Trace: src/VX_mem_coalescer.sv:112:5
	wire [((OUT_REQS * DATA_RATIO) * DATA_IN_WIDTH) - 1:0] req_data_merged;
	// Trace: src/VX_mem_coalescer.sv:113:5
	genvar _gv_i_70;
	generate
		for (_gv_i_70 = 0; _gv_i_70 < OUT_REQS; _gv_i_70 = _gv_i_70 + 1) begin : g_data_merged
			localparam i = _gv_i_70;
			// Trace: src/VX_mem_coalescer.sv:114:9
			reg [(DATA_RATIO * DATA_IN_SIZE) - 1:0] byteen_merged;
			// Trace: src/VX_mem_coalescer.sv:115:9
			reg [(DATA_RATIO * DATA_IN_WIDTH) - 1:0] data_merged;
			// Trace: src/VX_mem_coalescer.sv:116:9
			always @(*) begin
				// Trace: src/VX_mem_coalescer.sv:117:13
				byteen_merged = 1'sb0;
				// Trace: src/VX_mem_coalescer.sv:118:13
				data_merged = 1'sbx;
				// Trace: src/VX_mem_coalescer.sv:119:13
				begin : sv2v_autoblock_1
					// Trace: src/VX_mem_coalescer.sv:119:18
					integer j;
					// Trace: src/VX_mem_coalescer.sv:119:18
					for (j = 0; j < DATA_RATIO; j = j + 1)
						begin
							// Trace: src/VX_mem_coalescer.sv:120:17
							begin : sv2v_autoblock_2
								// Trace: src/VX_mem_coalescer.sv:120:22
								integer k;
								// Trace: src/VX_mem_coalescer.sv:120:22
								for (k = 0; k < DATA_IN_SIZE; k = k + 1)
									begin
										// Trace: src/VX_mem_coalescer.sv:121:21
										if (current_pmask[(i * DATA_RATIO) + j] && in_req_byteen[(((DATA_RATIO * i) + j) * DATA_IN_SIZE) + k]) begin
											// Trace: src/VX_mem_coalescer.sv:122:25
											byteen_merged[(in_addr_offset[((DATA_RATIO * i) + j) * DATA_RATIO_W+:DATA_RATIO_W] * DATA_IN_SIZE) + k] = 1'b1;
											// Trace: src/VX_mem_coalescer.sv:123:25
											data_merged[(in_addr_offset[((DATA_RATIO * i) + j) * DATA_RATIO_W+:DATA_RATIO_W] * DATA_IN_WIDTH) + (k * 8)+:8] = in_req_data[(((DATA_RATIO * i) + j) * DATA_IN_WIDTH) + (k * 8)+:8];
										end
									end
							end
						end
				end
			end
			// Trace: src/VX_mem_coalescer.sv:128:9
			assign req_byteen_merged[DATA_IN_SIZE * (i * DATA_RATIO)+:DATA_IN_SIZE * DATA_RATIO] = byteen_merged;
			// Trace: src/VX_mem_coalescer.sv:129:9
			assign req_data_merged[DATA_IN_WIDTH * (i * DATA_RATIO)+:DATA_IN_WIDTH * DATA_RATIO] = data_merged;
		end
	endgenerate
	// Trace: src/VX_mem_coalescer.sv:131:5
	wire is_last_batch = ~(|((in_req_mask & ~addr_matches_r) & req_rem_mask_r));
	// Trace: src/VX_mem_coalescer.sv:132:5
	wire out_req_fire = out_req_valid && out_req_ready;
	// Trace: src/VX_mem_coalescer.sv:133:5
	always @(*) begin
		// Trace: src/VX_mem_coalescer.sv:134:9
		state_n = state_r;
		// Trace: src/VX_mem_coalescer.sv:135:9
		out_req_valid_n = out_req_valid_r;
		// Trace: src/VX_mem_coalescer.sv:136:9
		out_req_mask_n = out_req_mask_r;
		// Trace: src/VX_mem_coalescer.sv:137:9
		out_req_rw_n = out_req_rw_r;
		// Trace: src/VX_mem_coalescer.sv:138:9
		out_req_addr_n = out_req_addr_r;
		// Trace: src/VX_mem_coalescer.sv:139:9
		out_req_flags_n = out_req_flags_r;
		// Trace: src/VX_mem_coalescer.sv:140:9
		out_req_byteen_n = out_req_byteen_r;
		// Trace: src/VX_mem_coalescer.sv:141:9
		out_req_data_n = out_req_data_r;
		// Trace: src/VX_mem_coalescer.sv:142:9
		out_req_tag_n = out_req_tag_r;
		// Trace: src/VX_mem_coalescer.sv:143:9
		req_rem_mask_n = req_rem_mask_r;
		// Trace: src/VX_mem_coalescer.sv:144:9
		in_req_ready_n = 0;
		// Trace: src/VX_mem_coalescer.sv:145:9
		case (state_r)
			STATE_WAIT: begin
				// Trace: src/VX_mem_coalescer.sv:147:13
				if (out_req_fire)
					// Trace: src/VX_mem_coalescer.sv:148:17
					out_req_valid_n = 0;
				if ((in_req_valid && ~out_req_valid_n) && ~ibuf_full)
					// Trace: src/VX_mem_coalescer.sv:151:17
					state_n = STATE_SEND;
			end
			default: begin
				// Trace: src/VX_mem_coalescer.sv:155:13
				state_n = STATE_WAIT;
				// Trace: src/VX_mem_coalescer.sv:156:13
				out_req_valid_n = 1;
				// Trace: src/VX_mem_coalescer.sv:157:13
				out_req_mask_n = batch_valid_r;
				// Trace: src/VX_mem_coalescer.sv:158:13
				out_req_rw_n = in_req_rw;
				// Trace: src/VX_mem_coalescer.sv:159:13
				out_req_addr_n = seed_addr_r;
				// Trace: src/VX_mem_coalescer.sv:160:13
				out_req_flags_n = seed_flags_r;
				// Trace: src/VX_mem_coalescer.sv:161:13
				out_req_byteen_n = req_byteen_merged;
				// Trace: src/VX_mem_coalescer.sv:162:13
				out_req_data_n = req_data_merged;
				// Trace: src/VX_mem_coalescer.sv:163:13
				out_req_tag_n = {in_req_tag[TAG_WIDTH - 1-:UUID_WIDTH], ibuf_waddr};
				// Trace: src/VX_mem_coalescer.sv:164:13
				req_rem_mask_n = (is_last_batch ? {NUM_REQS {1'sb1}} : req_rem_mask_r & ~current_pmask);
				// Trace: src/VX_mem_coalescer.sv:165:13
				in_req_ready_n = is_last_batch;
			end
		endcase
	end
	// Trace: src/VX_mem_coalescer.sv:169:5
	VX_pipe_register #(
		.DATAW(((((1 + NUM_REQS) + 2) + NUM_REQS) + (OUT_REQS * ((((((2 + OUT_ADDR_WIDTH) + (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) + OUT_ADDR_WIDTH) + (FLAGS_WIDTH > 0 ? FLAGS_WIDTH : 1)) + DATA_OUT_SIZE) + DATA_OUT_WIDTH))) + OUT_TAG_WIDTH),
		.RESETW((1 + NUM_REQS) + 1),
		.INIT_VALUE({1'b0, {NUM_REQS {1'b1}}, 1'b0})
	) pipe_reg(
		.clk(clk),
		.reset(reset),
		.enable(1'b1),
		.data_in({state_n, req_rem_mask_n, out_req_valid_n, out_req_rw_n, addr_matches_n, batch_valid_n, out_req_mask_n, seed_addr_n, seed_flags_n, out_req_addr_n, out_req_flags_n, out_req_byteen_n, out_req_data_n, out_req_tag_n}),
		.data_out({state_r, req_rem_mask_r, out_req_valid_r, out_req_rw_r, addr_matches_r, batch_valid_r, out_req_mask_r, seed_addr_r, seed_flags_r, out_req_addr_r, out_req_flags_r, out_req_byteen_r, out_req_data_r, out_req_tag_r})
	);
	// Trace: src/VX_mem_coalescer.sv:180:5
	wire out_rsp_fire = out_rsp_valid && out_rsp_ready;
	// Trace: src/VX_mem_coalescer.sv:181:5
	wire out_rsp_eop;
	// Trace: src/VX_mem_coalescer.sv:182:5
	wire req_sent = state_r == STATE_SEND;
	// Trace: src/VX_mem_coalescer.sv:183:5
	assign ibuf_push = req_sent && ~in_req_rw;
	// Trace: src/VX_mem_coalescer.sv:184:5
	assign ibuf_pop = out_rsp_fire && out_rsp_eop;
	// Trace: src/VX_mem_coalescer.sv:185:5
	assign ibuf_raddr = out_rsp_tag[QUEUE_ADDRW - 1:0];
	// Trace: src/VX_mem_coalescer.sv:186:5
	wire [TAG_ID_WIDTH - 1:0] ibuf_din_tag = in_req_tag[TAG_ID_WIDTH - 1:0];
	// Trace: src/VX_mem_coalescer.sv:187:5
	wire [(NUM_REQS * DATA_RATIO_W) - 1:0] ibuf_din_offset = in_addr_offset;
	// Trace: src/VX_mem_coalescer.sv:188:5
	wire [NUM_REQS - 1:0] ibuf_din_pmask = current_pmask;
	// Trace: src/VX_mem_coalescer.sv:189:5
	assign ibuf_din = {ibuf_din_tag, ibuf_din_pmask, ibuf_din_offset};
	// Trace: src/VX_mem_coalescer.sv:190:5
	VX_index_buffer #(
		.DATAW(IBUF_DATA_WIDTH),
		.SIZE(QUEUE_SIZE)
	) req_ibuf(
		.clk(clk),
		.reset(reset),
		.acquire_en(ibuf_push),
		.write_addr(ibuf_waddr),
		.write_data(ibuf_din),
		.read_data(ibuf_dout),
		.read_addr(ibuf_raddr),
		.release_en(ibuf_pop),
		.full(ibuf_full),
		.empty(ibuf_empty)
	);
	// Trace: src/VX_mem_coalescer.sv:205:5
	assign out_req_valid = out_req_valid_r;
	// Trace: src/VX_mem_coalescer.sv:206:5
	assign out_req_rw = out_req_rw_r;
	// Trace: src/VX_mem_coalescer.sv:207:5
	assign out_req_mask = out_req_mask_r;
	// Trace: src/VX_mem_coalescer.sv:208:5
	assign out_req_byteen = out_req_byteen_r;
	// Trace: src/VX_mem_coalescer.sv:209:5
	assign out_req_addr = out_req_addr_r;
	// Trace: src/VX_mem_coalescer.sv:210:5
	generate
		if (FLAGS_WIDTH != 0) begin : g_out_req_flags
			// Trace: src/VX_mem_coalescer.sv:211:9
			assign out_req_flags = out_req_flags_r;
		end
		else begin : g_out_req_flags_0
			// Trace: src/VX_mem_coalescer.sv:213:9
			assign out_req_flags = 1'sb0;
		end
	endgenerate
	// Trace: src/VX_mem_coalescer.sv:215:5
	assign out_req_data = out_req_data_r;
	// Trace: src/VX_mem_coalescer.sv:216:5
	assign out_req_tag = out_req_tag_r;
	// Trace: src/VX_mem_coalescer.sv:217:5
	assign in_req_ready = in_req_ready_n;
	// Trace: src/VX_mem_coalescer.sv:218:5
	reg [(QUEUE_SIZE * OUT_REQS) - 1:0] rsp_rem_mask;
	// Trace: src/VX_mem_coalescer.sv:219:5
	wire [OUT_REQS - 1:0] rsp_rem_mask_n = rsp_rem_mask[ibuf_raddr * OUT_REQS+:OUT_REQS] & ~out_rsp_mask;
	// Trace: src/VX_mem_coalescer.sv:220:5
	assign out_rsp_eop = ~(|rsp_rem_mask_n);
	// Trace: src/VX_mem_coalescer.sv:221:5
	always @(posedge clk) begin
		// Trace: src/VX_mem_coalescer.sv:222:9
		if (ibuf_push)
			// Trace: src/VX_mem_coalescer.sv:223:13
			rsp_rem_mask[ibuf_waddr * OUT_REQS+:OUT_REQS] <= batch_valid_r;
		if (out_rsp_fire)
			// Trace: src/VX_mem_coalescer.sv:226:13
			rsp_rem_mask[ibuf_raddr * OUT_REQS+:OUT_REQS] <= rsp_rem_mask_n;
	end
	// Trace: src/VX_mem_coalescer.sv:229:5
	wire [(NUM_REQS * DATA_RATIO_W) - 1:0] ibuf_dout_offset;
	// Trace: src/VX_mem_coalescer.sv:230:5
	wire [NUM_REQS - 1:0] ibuf_dout_pmask;
	// Trace: src/VX_mem_coalescer.sv:231:5
	wire [TAG_ID_WIDTH - 1:0] ibuf_dout_tag;
	// Trace: src/VX_mem_coalescer.sv:232:5
	assign {ibuf_dout_tag, ibuf_dout_pmask, ibuf_dout_offset} = ibuf_dout;
	// Trace: src/VX_mem_coalescer.sv:233:5
	wire [(NUM_REQS * DATA_IN_WIDTH) - 1:0] in_rsp_data_n;
	// Trace: src/VX_mem_coalescer.sv:234:5
	genvar _gv_i_71;
	generate
		for (_gv_i_71 = 0; _gv_i_71 < OUT_REQS; _gv_i_71 = _gv_i_71 + 1) begin : g_in_rsp_data_n
			localparam i = _gv_i_71;
			genvar _gv_j_10;
			for (_gv_j_10 = 0; _gv_j_10 < DATA_RATIO; _gv_j_10 = _gv_j_10 + 1) begin : g_j
				localparam j = _gv_j_10;
				// Trace: src/VX_mem_coalescer.sv:236:13
				assign in_rsp_data_n[((i * DATA_RATIO) + j) * DATA_IN_WIDTH+:DATA_IN_WIDTH] = out_rsp_data[(i * DATA_OUT_WIDTH) + (ibuf_dout_offset[((i * DATA_RATIO) + j) * DATA_RATIO_W+:DATA_RATIO_W] * DATA_IN_WIDTH)+:DATA_IN_WIDTH];
			end
		end
	endgenerate
	// Trace: src/VX_mem_coalescer.sv:239:5
	wire [NUM_REQS - 1:0] in_rsp_mask_n;
	// Trace: src/VX_mem_coalescer.sv:240:5
	genvar _gv_i_72;
	generate
		for (_gv_i_72 = 0; _gv_i_72 < OUT_REQS; _gv_i_72 = _gv_i_72 + 1) begin : g_in_rsp_mask_n
			localparam i = _gv_i_72;
			genvar _gv_j_11;
			for (_gv_j_11 = 0; _gv_j_11 < DATA_RATIO; _gv_j_11 = _gv_j_11 + 1) begin : g_j
				localparam j = _gv_j_11;
				// Trace: src/VX_mem_coalescer.sv:242:13
				assign in_rsp_mask_n[(i * DATA_RATIO) + j] = out_rsp_mask[i] && ibuf_dout_pmask[(i * DATA_RATIO) + j];
			end
		end
	endgenerate
	// Trace: src/VX_mem_coalescer.sv:245:5
	assign in_rsp_valid = out_rsp_valid;
	// Trace: src/VX_mem_coalescer.sv:246:5
	assign in_rsp_mask = in_rsp_mask_n;
	// Trace: src/VX_mem_coalescer.sv:247:5
	assign in_rsp_data = in_rsp_data_n;
	// Trace: src/VX_mem_coalescer.sv:248:5
	assign in_rsp_tag = {out_rsp_tag[OUT_TAG_WIDTH - 1-:UUID_WIDTH], ibuf_dout_tag};
	// Trace: src/VX_mem_coalescer.sv:249:5
	assign out_rsp_ready = in_rsp_ready;
	// Trace: src/VX_mem_coalescer.sv:250:5
	reg [PERF_CTR_BITS - 1:0] misses_r;
	// Trace: src/VX_mem_coalescer.sv:251:5
	wire partial_transfer = out_req_fire && (req_rem_mask_r != {NUM_REQS {1'sb1}});
	// Trace: src/VX_mem_coalescer.sv:252:5
	function automatic [PERF_CTR_BITS - 1:0] sv2v_cast_8BEE5;
		input reg [PERF_CTR_BITS - 1:0] inp;
		sv2v_cast_8BEE5 = inp;
	endfunction
	always @(posedge clk)
		// Trace: src/VX_mem_coalescer.sv:253:9
		if (reset)
			// Trace: src/VX_mem_coalescer.sv:254:13
			misses_r <= 1'sb0;
		else
			// Trace: src/VX_mem_coalescer.sv:256:13
			misses_r <= misses_r + sv2v_cast_8BEE5(partial_transfer);
	// Trace: src/VX_mem_coalescer.sv:259:5
	assign misses = misses_r;
endmodule
module VX_cache_flush (
	clk,
	reset,
	flush_begin,
	flush_end,
	flush_init,
	flush_valid,
	flush_line,
	flush_way,
	flush_ready,
	mshr_empty,
	bank_empty
);
	// removed import VX_gpu_pkg::*;
	// Trace: src/VX_cache_flush.sv:2:15
	parameter BANK_ID = 0;
	// Trace: src/VX_cache_flush.sv:3:15
	parameter CACHE_SIZE = 1024;
	// Trace: src/VX_cache_flush.sv:4:15
	parameter LINE_SIZE = 64;
	// Trace: src/VX_cache_flush.sv:5:15
	parameter NUM_BANKS = 1;
	// Trace: src/VX_cache_flush.sv:6:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_flush.sv:7:15
	parameter WRITEBACK = 0;
	// Trace: src/VX_cache_flush.sv:9:5
	input wire clk;
	// Trace: src/VX_cache_flush.sv:10:5
	input wire reset;
	// Trace: src/VX_cache_flush.sv:11:5
	input wire flush_begin;
	// Trace: src/VX_cache_flush.sv:12:5
	output wire flush_end;
	// Trace: src/VX_cache_flush.sv:13:5
	output wire flush_init;
	// Trace: src/VX_cache_flush.sv:14:5
	output wire flush_valid;
	// Trace: src/VX_cache_flush.sv:15:5
	output wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] flush_line;
	// Trace: src/VX_cache_flush.sv:16:5
	output wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] flush_way;
	// Trace: src/VX_cache_flush.sv:17:5
	input wire flush_ready;
	// Trace: src/VX_cache_flush.sv:18:5
	input wire mshr_empty;
	// Trace: src/VX_cache_flush.sv:19:5
	input wire bank_empty;
	// Trace: src/VX_cache_flush.sv:21:5
	localparam CTR_WIDTH = $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) + (WRITEBACK ? $clog2(NUM_WAYS) : 0);
	// Trace: src/VX_cache_flush.sv:22:5
	localparam STATE_IDLE = 0;
	// Trace: src/VX_cache_flush.sv:23:5
	localparam STATE_INIT = 1;
	// Trace: src/VX_cache_flush.sv:24:5
	localparam STATE_WAIT1 = 2;
	// Trace: src/VX_cache_flush.sv:25:5
	localparam STATE_FLUSH = 3;
	// Trace: src/VX_cache_flush.sv:26:5
	localparam STATE_WAIT2 = 4;
	// Trace: src/VX_cache_flush.sv:27:5
	localparam STATE_DONE = 5;
	// Trace: src/VX_cache_flush.sv:28:5
	reg [2:0] state;
	reg [2:0] state_n;
	// Trace: src/VX_cache_flush.sv:29:5
	reg [CTR_WIDTH - 1:0] counter;
	// Trace: src/VX_cache_flush.sv:30:5
	always @(*) begin
		// Trace: src/VX_cache_flush.sv:31:9
		state_n = state;
		// Trace: src/VX_cache_flush.sv:32:9
		case (state)
			default:
				// Trace: src/VX_cache_flush.sv:34:17
				if (flush_begin)
					// Trace: src/VX_cache_flush.sv:35:21
					state_n = STATE_WAIT1;
			STATE_INIT:
				// Trace: src/VX_cache_flush.sv:39:17
				if (counter == ((2 ** $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))
					// Trace: src/VX_cache_flush.sv:40:21
					state_n = STATE_IDLE;
			STATE_WAIT1:
				// Trace: src/VX_cache_flush.sv:44:17
				if (mshr_empty)
					// Trace: src/VX_cache_flush.sv:45:21
					state_n = STATE_FLUSH;
			STATE_FLUSH:
				// Trace: src/VX_cache_flush.sv:49:17
				if ((counter == ((2 ** CTR_WIDTH) - 1)) && flush_ready)
					// Trace: src/VX_cache_flush.sv:50:21
					state_n = (BANK_ID == 0 ? STATE_DONE : STATE_WAIT2);
			STATE_WAIT2:
				// Trace: src/VX_cache_flush.sv:54:17
				if (bank_empty)
					// Trace: src/VX_cache_flush.sv:55:21
					state_n = STATE_DONE;
			STATE_DONE:
				// Trace: src/VX_cache_flush.sv:59:17
				state_n = STATE_IDLE;
		endcase
	end
	// Trace: src/VX_cache_flush.sv:63:5
	function automatic signed [CTR_WIDTH - 1:0] sv2v_cast_8E811_signed;
		input reg signed [CTR_WIDTH - 1:0] inp;
		sv2v_cast_8E811_signed = inp;
	endfunction
	always @(posedge clk)
		// Trace: src/VX_cache_flush.sv:64:9
		if (reset) begin
			// Trace: src/VX_cache_flush.sv:65:13
			state <= STATE_INIT;
			// Trace: src/VX_cache_flush.sv:66:13
			counter <= 1'sb0;
		end
		else begin
			// Trace: src/VX_cache_flush.sv:68:13
			state <= state_n;
			// Trace: src/VX_cache_flush.sv:69:13
			if (state != STATE_IDLE) begin
				begin
					// Trace: src/VX_cache_flush.sv:70:17
					if ((state == STATE_INIT) || ((state == STATE_FLUSH) && flush_ready))
						// Trace: src/VX_cache_flush.sv:72:21
						counter <= counter + sv2v_cast_8E811_signed(1);
				end
			end
			else
				// Trace: src/VX_cache_flush.sv:75:17
				counter <= 1'sb0;
		end
	// Trace: src/VX_cache_flush.sv:79:5
	assign flush_end = state == STATE_DONE;
	// Trace: src/VX_cache_flush.sv:80:5
	assign flush_init = state == STATE_INIT;
	// Trace: src/VX_cache_flush.sv:81:5
	assign flush_valid = state == STATE_FLUSH;
	// Trace: src/VX_cache_flush.sv:82:5
	assign flush_line = counter[$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0];
	// Trace: src/VX_cache_flush.sv:83:5
	generate
		if (WRITEBACK && (NUM_WAYS > 1)) begin : g_flush_way
			// Trace: src/VX_cache_flush.sv:84:9
			assign flush_way = counter[$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))+:$clog2(NUM_WAYS)];
		end
		else begin : g_flush_way_all
			// Trace: src/VX_cache_flush.sv:86:9
			assign flush_way = 1'sb0;
		end
	endgenerate
endmodule
// removed module with interface ports: VX_fpu_unit
// removed module with interface ports: VX_execute
module VX_elastic_buffer (
	clk,
	reset,
	valid_in,
	ready_in,
	data_in,
	data_out,
	ready_out,
	valid_out
);
	// Trace: src/VX_elastic_buffer.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_elastic_buffer.sv:3:15
	parameter SIZE = 1;
	// Trace: src/VX_elastic_buffer.sv:4:15
	parameter OUT_REG = 0;
	// Trace: src/VX_elastic_buffer.sv:5:15
	parameter LUTRAM = 0;
	// Trace: src/VX_elastic_buffer.sv:7:5
	input wire clk;
	// Trace: src/VX_elastic_buffer.sv:8:5
	input wire reset;
	// Trace: src/VX_elastic_buffer.sv:9:5
	input wire valid_in;
	// Trace: src/VX_elastic_buffer.sv:10:5
	output wire ready_in;
	// Trace: src/VX_elastic_buffer.sv:11:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_elastic_buffer.sv:12:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_elastic_buffer.sv:13:5
	input wire ready_out;
	// Trace: src/VX_elastic_buffer.sv:14:5
	output wire valid_out;
	// Trace: src/VX_elastic_buffer.sv:16:5
	generate
		if (SIZE == 0) begin : g_passthru
			// Trace: src/VX_elastic_buffer.sv:17:9
			assign valid_out = valid_in;
			// Trace: src/VX_elastic_buffer.sv:18:9
			assign data_out = data_in;
			// Trace: src/VX_elastic_buffer.sv:19:9
			assign ready_in = ready_out;
		end
		else if (SIZE == 1) begin : g_eb1
			// Trace: src/VX_elastic_buffer.sv:21:9
			VX_pipe_buffer #(
				.DATAW(DATAW),
				.DEPTH((OUT_REG > 1 ? OUT_REG : 1))
			) pipe_buffer(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_in),
				.data_in(data_in),
				.ready_in(ready_in),
				.valid_out(valid_out),
				.data_out(data_out),
				.ready_out(ready_out)
			);
		end
		else if ((SIZE == 2) && (LUTRAM == 0)) begin : g_eb2
			// Trace: src/VX_elastic_buffer.sv:35:9
			wire valid_out_t;
			// Trace: src/VX_elastic_buffer.sv:36:9
			wire [DATAW - 1:0] data_out_t;
			// Trace: src/VX_elastic_buffer.sv:37:9
			wire ready_out_t;
			// Trace: src/VX_elastic_buffer.sv:38:9
			VX_stream_buffer #(
				.DATAW(DATAW),
				.OUT_REG(OUT_REG == 1)
			) stream_buffer(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_in),
				.data_in(data_in),
				.ready_in(ready_in),
				.valid_out(valid_out_t),
				.data_out(data_out_t),
				.ready_out(ready_out_t)
			);
			// Trace: src/VX_elastic_buffer.sv:51:9
			VX_pipe_buffer #(
				.DATAW(DATAW),
				.DEPTH((OUT_REG > 1 ? OUT_REG - 1 : 0))
			) out_buf(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_out_t),
				.data_in(data_out_t),
				.ready_in(ready_out_t),
				.valid_out(valid_out),
				.data_out(data_out),
				.ready_out(ready_out)
			);
		end
		else begin : g_ebN
			// Trace: src/VX_elastic_buffer.sv:65:9
			wire empty;
			wire full;
			// Trace: src/VX_elastic_buffer.sv:66:9
			wire [DATAW - 1:0] data_out_t;
			// Trace: src/VX_elastic_buffer.sv:67:9
			wire ready_out_t;
			// Trace: src/VX_elastic_buffer.sv:68:9
			wire valid_out_t = ~empty;
			// Trace: src/VX_elastic_buffer.sv:69:9
			wire push = valid_in && ready_in;
			// Trace: src/VX_elastic_buffer.sv:70:9
			wire pop = valid_out_t && ready_out_t;
			// Trace: src/VX_elastic_buffer.sv:71:9
			VX_fifo_queue #(
				.DATAW(DATAW),
				.DEPTH(SIZE),
				.OUT_REG(OUT_REG == 1),
				.LUTRAM(LUTRAM)
			) fifo_queue(
				.clk(clk),
				.reset(reset),
				.push(push),
				.pop(pop),
				.data_in(data_in),
				.data_out(data_out_t),
				.empty(empty),
				.full(full),
				.alm_empty(),
				.alm_full(),
				.size()
			);
			// Trace: src/VX_elastic_buffer.sv:89:9
			assign ready_in = ~full;
			// Trace: src/VX_elastic_buffer.sv:90:9
			VX_pipe_buffer #(
				.DATAW(DATAW),
				.DEPTH((OUT_REG > 1 ? OUT_REG - 1 : 0))
			) out_buf(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_out_t),
				.data_in(data_out_t),
				.ready_in(ready_out_t),
				.valid_out(valid_out),
				.data_out(data_out),
				.ready_out(ready_out)
			);
		end
	endgenerate
endmodule
module VX_cache_data (
	clk,
	reset,
	init,
	fill,
	flush,
	read,
	write,
	line_idx,
	evict_way,
	tag_matches,
	fill_data,
	write_word,
	write_byteen,
	word_idx,
	way_idx_r,
	read_data,
	evict_byteen
);
	// removed import VX_gpu_pkg::*;
	// Trace: src/VX_cache_data.sv:2:15
	parameter CACHE_SIZE = 1024;
	// Trace: src/VX_cache_data.sv:3:15
	parameter LINE_SIZE = 16;
	// Trace: src/VX_cache_data.sv:4:15
	parameter NUM_BANKS = 1;
	// Trace: src/VX_cache_data.sv:5:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_data.sv:6:15
	parameter WORD_SIZE = 1;
	// Trace: src/VX_cache_data.sv:7:15
	parameter WRITE_ENABLE = 1;
	// Trace: src/VX_cache_data.sv:8:15
	parameter WRITEBACK = 0;
	// Trace: src/VX_cache_data.sv:9:15
	parameter DIRTY_BYTES = 0;
	// Trace: src/VX_cache_data.sv:11:5
	input wire clk;
	// Trace: src/VX_cache_data.sv:12:5
	input wire reset;
	// Trace: src/VX_cache_data.sv:13:5
	input wire init;
	// Trace: src/VX_cache_data.sv:14:5
	input wire fill;
	// Trace: src/VX_cache_data.sv:15:5
	input wire flush;
	// Trace: src/VX_cache_data.sv:16:5
	input wire read;
	// Trace: src/VX_cache_data.sv:17:5
	input wire write;
	// Trace: src/VX_cache_data.sv:18:5
	input wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] line_idx;
	// Trace: src/VX_cache_data.sv:19:5
	input wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] evict_way;
	// Trace: src/VX_cache_data.sv:20:5
	input wire [NUM_WAYS - 1:0] tag_matches;
	// Trace: src/VX_cache_data.sv:21:5
	input wire [((LINE_SIZE / WORD_SIZE) * (8 * WORD_SIZE)) - 1:0] fill_data;
	// Trace: src/VX_cache_data.sv:22:5
	input wire [(8 * WORD_SIZE) - 1:0] write_word;
	// Trace: src/VX_cache_data.sv:23:5
	input wire [WORD_SIZE - 1:0] write_byteen;
	// Trace: src/VX_cache_data.sv:24:5
	input wire [($clog2(LINE_SIZE / WORD_SIZE) > 0 ? $clog2(LINE_SIZE / WORD_SIZE) : 1) - 1:0] word_idx;
	// Trace: src/VX_cache_data.sv:25:5
	input wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] way_idx_r;
	// Trace: src/VX_cache_data.sv:26:5
	output wire [(8 * LINE_SIZE) - 1:0] read_data;
	// Trace: src/VX_cache_data.sv:27:5
	output wire [LINE_SIZE - 1:0] evict_byteen;
	// Trace: src/VX_cache_data.sv:29:5
	wire [((LINE_SIZE / WORD_SIZE) * WORD_SIZE) - 1:0] write_mask;
	// Trace: src/VX_cache_data.sv:30:5
	genvar _gv_i_73;
	generate
		for (_gv_i_73 = 0; _gv_i_73 < (LINE_SIZE / WORD_SIZE); _gv_i_73 = _gv_i_73 + 1) begin : g_write_mask
			localparam i = _gv_i_73;
			// Trace: src/VX_cache_data.sv:31:9
			wire word_en = ((LINE_SIZE / WORD_SIZE) == 1) || (word_idx == i);
			// Trace: src/VX_cache_data.sv:32:9
			assign write_mask[i * WORD_SIZE+:WORD_SIZE] = write_byteen & {WORD_SIZE {word_en}};
		end
	endgenerate
	// Trace: src/VX_cache_data.sv:34:5
	generate
		if (DIRTY_BYTES != 0) begin : g_dirty_bytes
			// Trace: src/VX_cache_data.sv:35:9
			wire [(NUM_WAYS * LINE_SIZE) - 1:0] byteen_rdata;
			genvar _gv_i_74;
			for (_gv_i_74 = 0; _gv_i_74 < NUM_WAYS; _gv_i_74 = _gv_i_74 + 1) begin : g_byteen_store
				localparam i = _gv_i_74;
				// Trace: src/VX_cache_data.sv:37:13
				wire [LINE_SIZE - 1:0] byteen_wdata = {LINE_SIZE {write}};
				// Trace: src/VX_cache_data.sv:38:13
				wire [LINE_SIZE - 1:0] byteen_wren = {LINE_SIZE {(init || fill) || flush}} | write_mask;
				// Trace: src/VX_cache_data.sv:39:13
				wire byteen_write = (((fill || flush) && ((NUM_WAYS == 1) || (evict_way == i))) || (write && tag_matches[i])) || init;
				// Trace: src/VX_cache_data.sv:42:13
				wire byteen_read = fill || flush;
				// Trace: src/VX_cache_data.sv:43:13
				VX_sp_ram #(
					.DATAW(LINE_SIZE),
					.WRENW(LINE_SIZE),
					.SIZE((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)),
					.OUT_REG(1),
					.RDW_MODE("R")
				) byteen_store(
					.clk(clk),
					.reset(reset),
					.read(byteen_read),
					.write(byteen_write),
					.wren(byteen_wren),
					.addr(line_idx),
					.wdata(byteen_wdata),
					.rdata(byteen_rdata[i * LINE_SIZE+:LINE_SIZE])
				);
			end
			// Trace: src/VX_cache_data.sv:60:9
			assign evict_byteen = byteen_rdata[way_idx_r * LINE_SIZE+:LINE_SIZE];
		end
		else begin : g_no_dirty_bytes
			// Trace: src/VX_cache_data.sv:62:9
			assign evict_byteen = 1'sb1;
		end
	endgenerate
	// Trace: src/VX_cache_data.sv:64:5
	wire [((NUM_WAYS * (LINE_SIZE / WORD_SIZE)) * (8 * WORD_SIZE)) - 1:0] line_rdata;
	// Trace: src/VX_cache_data.sv:65:5
	genvar _gv_i_75;
	generate
		for (_gv_i_75 = 0; _gv_i_75 < NUM_WAYS; _gv_i_75 = _gv_i_75 + 1) begin : g_data_store
			localparam i = _gv_i_75;
			// Trace: src/VX_cache_data.sv:66:9
			localparam WRENW = (WRITE_ENABLE ? LINE_SIZE : 1);
			// Trace: src/VX_cache_data.sv:67:9
			wire [((LINE_SIZE / WORD_SIZE) * (8 * WORD_SIZE)) - 1:0] line_wdata;
			// Trace: src/VX_cache_data.sv:68:9
			wire [WRENW - 1:0] line_wren;
			if (WRITE_ENABLE) begin : g_wren
				// Trace: src/VX_cache_data.sv:70:13
				assign line_wdata = (fill ? fill_data : {LINE_SIZE / WORD_SIZE {write_word}});
				// Trace: src/VX_cache_data.sv:71:13
				assign line_wren = {LINE_SIZE {fill}} | write_mask;
			end
			else begin : g_no_wren
				// Trace: src/VX_cache_data.sv:73:13
				assign line_wdata = fill_data;
				// Trace: src/VX_cache_data.sv:74:13
				assign line_wren = 1'b1;
			end
			// Trace: src/VX_cache_data.sv:76:9
			wire line_write = (fill && ((NUM_WAYS == 1) || (evict_way == i))) || ((write && tag_matches[i]) && WRITE_ENABLE);
			// Trace: src/VX_cache_data.sv:78:9
			wire line_read = read || ((fill || flush) && WRITEBACK);
			// Trace: src/VX_cache_data.sv:79:9
			VX_sp_ram #(
				.DATAW(8 * LINE_SIZE),
				.SIZE((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)),
				.WRENW(WRENW),
				.OUT_REG(1),
				.RDW_MODE("R")
			) data_store(
				.clk(clk),
				.reset(reset),
				.read(line_read),
				.write(line_write),
				.wren(line_wren),
				.addr(line_idx),
				.wdata(line_wdata),
				.rdata(line_rdata[(8 * WORD_SIZE) * (i * (LINE_SIZE / WORD_SIZE))+:(8 * WORD_SIZE) * (LINE_SIZE / WORD_SIZE)])
			);
		end
	endgenerate
	// Trace: src/VX_cache_data.sv:96:5
	assign read_data = line_rdata[(8 * WORD_SIZE) * (way_idx_r * (LINE_SIZE / WORD_SIZE))+:(8 * WORD_SIZE) * (LINE_SIZE / WORD_SIZE)];
endmodule
module VX_matrix_arbiter (
	clk,
	reset,
	requests,
	grant_index,
	grant_onehot,
	grant_valid,
	grant_ready
);
	// Trace: src/VX_matrix_arbiter.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_matrix_arbiter.sv:3:15
	parameter STICKY = 0;
	// Trace: src/VX_matrix_arbiter.sv:4:15
	parameter LOG_NUM_REQS = (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1);
	// Trace: src/VX_matrix_arbiter.sv:6:5
	input wire clk;
	// Trace: src/VX_matrix_arbiter.sv:7:5
	input wire reset;
	// Trace: src/VX_matrix_arbiter.sv:8:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: src/VX_matrix_arbiter.sv:9:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: src/VX_matrix_arbiter.sv:10:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: src/VX_matrix_arbiter.sv:11:5
	output wire grant_valid;
	// Trace: src/VX_matrix_arbiter.sv:12:5
	input wire grant_ready;
	// Trace: src/VX_matrix_arbiter.sv:14:5
	generate
		if (NUM_REQS == 1) begin : g_passthru
			// Trace: src/VX_matrix_arbiter.sv:15:9
			assign grant_index = 1'sb0;
			// Trace: src/VX_matrix_arbiter.sv:16:9
			assign grant_onehot = requests;
			// Trace: src/VX_matrix_arbiter.sv:17:9
			assign grant_valid = requests[0];
		end
		else begin : g_arbiter
			// Trace: src/VX_matrix_arbiter.sv:19:9
			reg [NUM_REQS - 1:1] state [NUM_REQS - 1:0];
			// Trace: src/VX_matrix_arbiter.sv:20:9
			wire [NUM_REQS - 1:0] pri [NUM_REQS - 1:0];
			// Trace: src/VX_matrix_arbiter.sv:21:9
			wire [NUM_REQS - 1:0] grant;
			// Trace: src/VX_matrix_arbiter.sv:22:9
			reg [NUM_REQS - 1:0] prev_grant;
			// Trace: src/VX_matrix_arbiter.sv:23:9
			always @(posedge clk)
				// Trace: src/VX_matrix_arbiter.sv:24:13
				if (reset)
					// Trace: src/VX_matrix_arbiter.sv:25:17
					prev_grant <= 1'sb0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_matrix_arbiter.sv:27:17
					prev_grant <= grant_onehot;
			// Trace: src/VX_matrix_arbiter.sv:30:9
			wire retain_grant = (STICKY != 0) && |(prev_grant & requests);
			// Trace: src/VX_matrix_arbiter.sv:31:9
			wire [NUM_REQS - 1:0] grant_w = (retain_grant ? prev_grant : grant);
			genvar _gv_r_4;
			for (_gv_r_4 = 0; _gv_r_4 < NUM_REQS; _gv_r_4 = _gv_r_4 + 1) begin : g_pri_r
				localparam r = _gv_r_4;
				genvar _gv_c_1;
				for (_gv_c_1 = 0; _gv_c_1 < NUM_REQS; _gv_c_1 = _gv_c_1 + 1) begin : g_pri_c
					localparam c = _gv_c_1;
					if (r > c) begin : g_row
						// Trace: src/VX_matrix_arbiter.sv:35:21
						assign pri[r][c] = requests[c] && state[c][r];
					end
					else if (r < c) begin : g_col
						// Trace: src/VX_matrix_arbiter.sv:37:21
						assign pri[r][c] = requests[c] && !state[r][c];
					end
					else begin : g_equal
						// Trace: src/VX_matrix_arbiter.sv:39:21
						assign pri[r][c] = 0;
					end
				end
			end
			genvar _gv_r_5;
			for (_gv_r_5 = 0; _gv_r_5 < NUM_REQS; _gv_r_5 = _gv_r_5 + 1) begin : g_grant
				localparam r = _gv_r_5;
				// Trace: src/VX_matrix_arbiter.sv:44:13
				assign grant[r] = requests[r] && ~(|pri[r]);
			end
			genvar _gv_r_6;
			for (_gv_r_6 = 0; _gv_r_6 < NUM_REQS; _gv_r_6 = _gv_r_6 + 1) begin : g_state_r
				localparam r = _gv_r_6;
				genvar _gv_c_2;
				for (_gv_c_2 = r + 1; _gv_c_2 < NUM_REQS; _gv_c_2 = _gv_c_2 + 1) begin : g_state_c
					localparam c = _gv_c_2;
					// Trace: src/VX_matrix_arbiter.sv:48:17
					always @(posedge clk)
						// Trace: src/VX_matrix_arbiter.sv:49:21
						if (reset)
							// Trace: src/VX_matrix_arbiter.sv:50:25
							state[r][c] <= 1'sb0;
						else if ((grant_valid && grant_ready) && ~retain_grant)
							// Trace: src/VX_matrix_arbiter.sv:52:25
							state[r][c] <= (state[r][c] || grant[c]) && ~grant[r];
				end
			end
			// Trace: src/VX_matrix_arbiter.sv:57:9
			assign grant_onehot = grant_w;
			// Trace: src/VX_matrix_arbiter.sv:58:9
			wire grant_valid_w;
			// Trace: src/VX_matrix_arbiter.sv:59:9
			VX_onehot_encoder #(.N(NUM_REQS)) encoder(
				.data_in(grant_w),
				.data_out(grant_index),
				.valid_out(grant_valid_w)
			);
			// Trace: src/VX_matrix_arbiter.sv:66:9
			assign grant_valid = (STICKY != 0 ? |requests : grant_valid_w);
		end
	endgenerate
endmodule
// removed module with interface ports: VX_alu_muldiv
// removed module with interface ports: VX_commit
module VX_stream_arb (
	clk,
	reset,
	valid_in,
	data_in,
	ready_in,
	valid_out,
	data_out,
	ready_out,
	sel_out
);
	// Trace: src/VX_stream_arb.sv:2:15
	parameter NUM_INPUTS = 1;
	// Trace: src/VX_stream_arb.sv:3:15
	parameter NUM_OUTPUTS = 1;
	// Trace: src/VX_stream_arb.sv:4:15
	parameter DATAW = 1;
	// Trace: src/VX_stream_arb.sv:5:15
	parameter STICKY = 0;
	// Trace: src/VX_stream_arb.sv:6:15
	parameter ARBITER = "R";
	// Trace: src/VX_stream_arb.sv:7:15
	parameter MAX_FANOUT = 8;
	// Trace: src/VX_stream_arb.sv:8:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_stream_arb.sv:9:15
	parameter NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? ((NUM_INPUTS + NUM_OUTPUTS) - 1) / NUM_OUTPUTS : ((NUM_OUTPUTS + NUM_INPUTS) - 1) / NUM_INPUTS);
	// Trace: src/VX_stream_arb.sv:10:15
	parameter SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
	// Trace: src/VX_stream_arb.sv:11:15
	parameter LOG_NUM_REQS = $clog2(NUM_REQS);
	// Trace: src/VX_stream_arb.sv:12:15
	parameter NUM_REQS_W = (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1);
	// Trace: src/VX_stream_arb.sv:14:5
	input wire clk;
	// Trace: src/VX_stream_arb.sv:15:5
	input wire reset;
	// Trace: src/VX_stream_arb.sv:16:5
	input wire [NUM_INPUTS - 1:0] valid_in;
	// Trace: src/VX_stream_arb.sv:17:5
	input wire [(NUM_INPUTS * DATAW) - 1:0] data_in;
	// Trace: src/VX_stream_arb.sv:18:5
	output wire [NUM_INPUTS - 1:0] ready_in;
	// Trace: src/VX_stream_arb.sv:19:5
	output wire [NUM_OUTPUTS - 1:0] valid_out;
	// Trace: src/VX_stream_arb.sv:20:5
	output wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out;
	// Trace: src/VX_stream_arb.sv:21:5
	input wire [NUM_OUTPUTS - 1:0] ready_out;
	// Trace: src/VX_stream_arb.sv:22:5
	output wire [(SEL_COUNT * NUM_REQS_W) - 1:0] sel_out;
	// Trace: src/VX_stream_arb.sv:24:5
	function automatic signed [NUM_REQS_W - 1:0] sv2v_cast_A9560_signed;
		input reg signed [NUM_REQS_W - 1:0] inp;
		sv2v_cast_A9560_signed = inp;
	endfunction
	generate
		if (NUM_INPUTS > NUM_OUTPUTS) begin : g_input_select
			if ((MAX_FANOUT != 0) && (NUM_REQS > (MAX_FANOUT + (MAX_FANOUT / 2)))) begin : g_fanout
				// Trace: src/VX_stream_arb.sv:26:13
				localparam NUM_SLICES = ((NUM_REQS + MAX_FANOUT) - 1) / MAX_FANOUT;
				// Trace: src/VX_stream_arb.sv:27:13
				localparam LOG_NUM_REQS2 = $clog2(MAX_FANOUT);
				// Trace: src/VX_stream_arb.sv:28:13
				localparam LOG_NUM_REQS3 = $clog2(NUM_SLICES);
				// Trace: src/VX_stream_arb.sv:29:13
				localparam DATAW2 = DATAW + LOG_NUM_REQS2;
				// Trace: src/VX_stream_arb.sv:30:13
				wire [(NUM_SLICES * NUM_OUTPUTS) - 1:0] valid_tmp;
				// Trace: src/VX_stream_arb.sv:31:13
				wire [((NUM_SLICES * NUM_OUTPUTS) * DATAW2) - 1:0] data_tmp;
				// Trace: src/VX_stream_arb.sv:32:13
				wire [(NUM_SLICES * NUM_OUTPUTS) - 1:0] ready_tmp;
				genvar _gv_s_2;
				for (_gv_s_2 = 0; _gv_s_2 < NUM_SLICES; _gv_s_2 = _gv_s_2 + 1) begin : g_slice_arbs
					localparam s = _gv_s_2;
					// Trace: src/VX_stream_arb.sv:34:17
					localparam SLICE_STRIDE = MAX_FANOUT * NUM_OUTPUTS;
					// Trace: src/VX_stream_arb.sv:35:17
					localparam SLICE_BEGIN = s * SLICE_STRIDE;
					// Trace: src/VX_stream_arb.sv:36:17
					localparam SLICE_END = ((SLICE_BEGIN + SLICE_STRIDE) < NUM_INPUTS ? SLICE_BEGIN + SLICE_STRIDE : NUM_INPUTS);
					// Trace: src/VX_stream_arb.sv:37:17
					localparam SLICE_SIZE = SLICE_END - SLICE_BEGIN;
					// Trace: src/VX_stream_arb.sv:38:17
					wire [(NUM_OUTPUTS * DATAW) - 1:0] data_tmp_u;
					// Trace: src/VX_stream_arb.sv:39:17
					wire [(NUM_OUTPUTS * LOG_NUM_REQS2) - 1:0] sel_tmp_u;
					// Trace: src/VX_stream_arb.sv:40:17
					VX_stream_arb #(
						.NUM_INPUTS(SLICE_SIZE),
						.NUM_OUTPUTS(NUM_OUTPUTS),
						.DATAW(DATAW),
						.ARBITER(ARBITER),
						.STICKY(STICKY),
						.MAX_FANOUT(MAX_FANOUT),
						.OUT_BUF(3)
					) fanout_slice_arb(
						.clk(clk),
						.reset(reset),
						.valid_in(valid_in[SLICE_END - 1:SLICE_BEGIN]),
						.data_in(data_in[DATAW * (((SLICE_END - 1) >= SLICE_BEGIN ? SLICE_END - 1 : ((SLICE_END - 1) + ((SLICE_END - 1) >= SLICE_BEGIN ? ((SLICE_END - 1) - SLICE_BEGIN) + 1 : (SLICE_BEGIN - (SLICE_END - 1)) + 1)) - 1) - (((SLICE_END - 1) >= SLICE_BEGIN ? ((SLICE_END - 1) - SLICE_BEGIN) + 1 : (SLICE_BEGIN - (SLICE_END - 1)) + 1) - 1))+:DATAW * ((SLICE_END - 1) >= SLICE_BEGIN ? ((SLICE_END - 1) - SLICE_BEGIN) + 1 : (SLICE_BEGIN - (SLICE_END - 1)) + 1)]),
						.ready_in(ready_in[SLICE_END - 1:SLICE_BEGIN]),
						.valid_out(valid_tmp[s * NUM_OUTPUTS+:NUM_OUTPUTS]),
						.data_out(data_tmp_u),
						.ready_out(ready_tmp[s * NUM_OUTPUTS+:NUM_OUTPUTS]),
						.sel_out(sel_tmp_u)
					);
					genvar _gv_o_1;
					for (_gv_o_1 = 0; _gv_o_1 < NUM_OUTPUTS; _gv_o_1 = _gv_o_1 + 1) begin : g_data_tmp
						localparam o = _gv_o_1;
						// Trace: src/VX_stream_arb.sv:60:21
						assign data_tmp[((s * NUM_OUTPUTS) + o) * DATAW2+:DATAW2] = {data_tmp_u[o * DATAW+:DATAW], sel_tmp_u[o * LOG_NUM_REQS2+:LOG_NUM_REQS2]};
					end
				end
				// Trace: src/VX_stream_arb.sv:63:13
				wire [(NUM_OUTPUTS * DATAW2) - 1:0] data_out_u;
				// Trace: src/VX_stream_arb.sv:64:13
				wire [(NUM_OUTPUTS * LOG_NUM_REQS3) - 1:0] sel_out_u;
				// Trace: src/VX_stream_arb.sv:65:13
				VX_stream_arb #(
					.NUM_INPUTS(NUM_SLICES * NUM_OUTPUTS),
					.NUM_OUTPUTS(NUM_OUTPUTS),
					.DATAW(DATAW2),
					.ARBITER(ARBITER),
					.STICKY(STICKY),
					.MAX_FANOUT(MAX_FANOUT),
					.OUT_BUF(OUT_BUF)
				) fanout_join_arb(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_tmp),
					.ready_in(ready_tmp),
					.data_in(data_tmp),
					.data_out(data_out_u),
					.sel_out(sel_out_u),
					.valid_out(valid_out),
					.ready_out(ready_out)
				);
				genvar _gv_o_2;
				for (_gv_o_2 = 0; _gv_o_2 < NUM_OUTPUTS; _gv_o_2 = _gv_o_2 + 1) begin : g_data_out
					localparam o = _gv_o_2;
					// Trace: src/VX_stream_arb.sv:85:17
					assign sel_out[o * NUM_REQS_W+:NUM_REQS_W] = {sel_out_u[o * LOG_NUM_REQS3+:LOG_NUM_REQS3], data_out_u[(o * DATAW2) + (LOG_NUM_REQS2 - 1)-:LOG_NUM_REQS2]};
					// Trace: src/VX_stream_arb.sv:86:17
					assign data_out[o * DATAW+:DATAW] = data_out_u[(o * DATAW2) + ((DATAW2 - 1) >= LOG_NUM_REQS2 ? DATAW2 - 1 : ((DATAW2 - 1) + ((DATAW2 - 1) >= LOG_NUM_REQS2 ? ((DATAW2 - 1) - LOG_NUM_REQS2) + 1 : (LOG_NUM_REQS2 - (DATAW2 - 1)) + 1)) - 1)-:((DATAW2 - 1) >= LOG_NUM_REQS2 ? ((DATAW2 - 1) - LOG_NUM_REQS2) + 1 : (LOG_NUM_REQS2 - (DATAW2 - 1)) + 1)];
				end
			end
			else begin : g_arbiter
				// Trace: src/VX_stream_arb.sv:89:13
				wire [NUM_REQS - 1:0] arb_requests;
				// Trace: src/VX_stream_arb.sv:90:13
				wire arb_valid;
				// Trace: src/VX_stream_arb.sv:91:13
				wire [NUM_REQS_W - 1:0] arb_index;
				// Trace: src/VX_stream_arb.sv:92:13
				wire [NUM_REQS - 1:0] arb_onehot;
				// Trace: src/VX_stream_arb.sv:93:13
				wire arb_ready;
				genvar _gv_r_7;
				for (_gv_r_7 = 0; _gv_r_7 < NUM_REQS; _gv_r_7 = _gv_r_7 + 1) begin : g_requests
					localparam r = _gv_r_7;
					// Trace: src/VX_stream_arb.sv:95:17
					wire [NUM_OUTPUTS - 1:0] requests;
					genvar _gv_o_3;
					for (_gv_o_3 = 0; _gv_o_3 < NUM_OUTPUTS; _gv_o_3 = _gv_o_3 + 1) begin : g_o
						localparam o = _gv_o_3;
						// Trace: src/VX_stream_arb.sv:97:21
						localparam i = (r * NUM_OUTPUTS) + o;
						// Trace: src/VX_stream_arb.sv:98:21
						assign requests[o] = valid_in[i];
					end
					// Trace: src/VX_stream_arb.sv:100:17
					assign arb_requests[r] = |requests;
				end
				// Trace: src/VX_stream_arb.sv:102:13
				VX_generic_arbiter #(
					.NUM_REQS(NUM_REQS),
					.TYPE(ARBITER),
					.STICKY(STICKY)
				) arbiter(
					.clk(clk),
					.reset(reset),
					.requests(arb_requests),
					.grant_valid(arb_valid),
					.grant_index(arb_index),
					.grant_onehot(arb_onehot),
					.grant_ready(arb_ready)
				);
				// Trace: src/VX_stream_arb.sv:115:13
				wire [NUM_OUTPUTS - 1:0] valid_out_w;
				// Trace: src/VX_stream_arb.sv:116:13
				wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out_w;
				// Trace: src/VX_stream_arb.sv:117:13
				wire [NUM_OUTPUTS - 1:0] ready_out_w;
				genvar _gv_o_4;
				for (_gv_o_4 = 0; _gv_o_4 < NUM_OUTPUTS; _gv_o_4 = _gv_o_4 + 1) begin : g_data_out_w
					localparam o = _gv_o_4;
					// Trace: src/VX_stream_arb.sv:119:17
					wire [NUM_REQS - 1:0] valid_in_w;
					// Trace: src/VX_stream_arb.sv:120:17
					wire [(NUM_REQS * DATAW) - 1:0] data_in_w;
					genvar _gv_r_8;
					for (_gv_r_8 = 0; _gv_r_8 < NUM_REQS; _gv_r_8 = _gv_r_8 + 1) begin : g_r
						localparam r = _gv_r_8;
						// Trace: src/VX_stream_arb.sv:122:21
						localparam i = (r * NUM_OUTPUTS) + o;
						if (r < NUM_INPUTS) begin : g_valid
							// Trace: src/VX_stream_arb.sv:124:25
							assign valid_in_w[r] = valid_in[i];
							// Trace: src/VX_stream_arb.sv:125:25
							assign data_in_w[r * DATAW+:DATAW] = data_in[i * DATAW+:DATAW];
						end
						else begin : g_padding
							// Trace: src/VX_stream_arb.sv:127:25
							assign valid_in_w[r] = 0;
							// Trace: src/VX_stream_arb.sv:128:25
							assign data_in_w[r * DATAW+:DATAW] = 1'sb0;
						end
					end
					// Trace: src/VX_stream_arb.sv:131:17
					assign valid_out_w[o] = (NUM_OUTPUTS == 1 ? arb_valid : |(valid_in_w & arb_onehot));
					// Trace: src/VX_stream_arb.sv:132:17
					assign data_out_w[o * DATAW+:DATAW] = data_in_w[arb_index * DATAW+:DATAW];
				end
				genvar _gv_i_84;
				for (_gv_i_84 = 0; _gv_i_84 < NUM_INPUTS; _gv_i_84 = _gv_i_84 + 1) begin : g_ready_in
					localparam i = _gv_i_84;
					// Trace: src/VX_stream_arb.sv:135:17
					localparam o = i % NUM_OUTPUTS;
					// Trace: src/VX_stream_arb.sv:136:17
					localparam r = i / NUM_OUTPUTS;
					// Trace: src/VX_stream_arb.sv:137:17
					assign ready_in[i] = ready_out_w[o] && arb_onehot[r];
				end
				// Trace: src/VX_stream_arb.sv:139:13
				assign arb_ready = |ready_out_w;
				genvar _gv_o_5;
				for (_gv_o_5 = 0; _gv_o_5 < NUM_OUTPUTS; _gv_o_5 = _gv_o_5 + 1) begin : g_out_buf
					localparam o = _gv_o_5;
					// Trace: src/VX_stream_arb.sv:141:17
					VX_elastic_buffer #(
						.DATAW(LOG_NUM_REQS + DATAW),
						.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
						.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2)),
						.LUTRAM((OUT_BUF & 8) != 0)
					) out_buf(
						.clk(clk),
						.reset(reset),
						.valid_in(valid_out_w[o]),
						.ready_in(ready_out_w[o]),
						.data_in({arb_index, data_out_w[o * DATAW+:DATAW]}),
						.data_out({sel_out[o * NUM_REQS_W+:NUM_REQS_W], data_out[o * DATAW+:DATAW]}),
						.valid_out(valid_out[o]),
						.ready_out(ready_out[o])
					);
				end
			end
		end
		else if (NUM_INPUTS < NUM_OUTPUTS) begin : g_output_select
			if ((MAX_FANOUT != 0) && (NUM_REQS > (MAX_FANOUT + (MAX_FANOUT / 2)))) begin : g_fanout
				// Trace: src/VX_stream_arb.sv:160:13
				localparam NUM_SLICES = ((NUM_REQS + MAX_FANOUT) - 1) / MAX_FANOUT;
				// Trace: src/VX_stream_arb.sv:161:13
				localparam LOG_NUM_REQS2 = $clog2(MAX_FANOUT);
				// Trace: src/VX_stream_arb.sv:162:13
				localparam LOG_NUM_REQS3 = $clog2(NUM_SLICES);
				// Trace: src/VX_stream_arb.sv:163:13
				wire [(NUM_SLICES * NUM_INPUTS) - 1:0] valid_tmp;
				// Trace: src/VX_stream_arb.sv:164:13
				wire [((NUM_SLICES * NUM_INPUTS) * DATAW) - 1:0] data_tmp;
				// Trace: src/VX_stream_arb.sv:165:13
				wire [(NUM_SLICES * NUM_INPUTS) - 1:0] ready_tmp;
				// Trace: src/VX_stream_arb.sv:166:13
				wire [(NUM_INPUTS * LOG_NUM_REQS3) - 1:0] sel_tmp;
				// Trace: src/VX_stream_arb.sv:167:13
				VX_stream_arb #(
					.NUM_INPUTS(NUM_INPUTS),
					.NUM_OUTPUTS(NUM_SLICES * NUM_INPUTS),
					.DATAW(DATAW),
					.ARBITER(ARBITER),
					.STICKY(STICKY),
					.MAX_FANOUT(MAX_FANOUT),
					.OUT_BUF(3)
				) fanout_fork_arb(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_in),
					.ready_in(ready_in),
					.data_in(data_in),
					.data_out(data_tmp),
					.valid_out(valid_tmp),
					.ready_out(ready_tmp),
					.sel_out(sel_tmp)
				);
				// Trace: src/VX_stream_arb.sv:186:13
				wire [((NUM_SLICES * NUM_INPUTS) * LOG_NUM_REQS2) - 1:0] sel_out_w;
				genvar _gv_s_3;
				for (_gv_s_3 = 0; _gv_s_3 < NUM_SLICES; _gv_s_3 = _gv_s_3 + 1) begin : g_slice_arbs
					localparam s = _gv_s_3;
					// Trace: src/VX_stream_arb.sv:188:17
					localparam SLICE_STRIDE = MAX_FANOUT * NUM_INPUTS;
					// Trace: src/VX_stream_arb.sv:189:17
					localparam SLICE_BEGIN = s * SLICE_STRIDE;
					// Trace: src/VX_stream_arb.sv:190:17
					localparam SLICE_END = ((SLICE_BEGIN + SLICE_STRIDE) < NUM_OUTPUTS ? SLICE_BEGIN + SLICE_STRIDE : NUM_OUTPUTS);
					// Trace: src/VX_stream_arb.sv:191:17
					localparam SLICE_SIZE = SLICE_END - SLICE_BEGIN;
					// Trace: src/VX_stream_arb.sv:192:17
					wire [(NUM_INPUTS * LOG_NUM_REQS2) - 1:0] sel_out_u;
					// Trace: src/VX_stream_arb.sv:193:17
					VX_stream_arb #(
						.NUM_INPUTS(NUM_INPUTS),
						.NUM_OUTPUTS(SLICE_SIZE),
						.DATAW(DATAW),
						.ARBITER(ARBITER),
						.STICKY(STICKY),
						.MAX_FANOUT(MAX_FANOUT),
						.OUT_BUF(OUT_BUF)
					) fanout_slice_arb(
						.clk(clk),
						.reset(reset),
						.valid_in(valid_tmp[s * NUM_INPUTS+:NUM_INPUTS]),
						.ready_in(ready_tmp[s * NUM_INPUTS+:NUM_INPUTS]),
						.data_in(data_tmp[DATAW * (s * NUM_INPUTS)+:DATAW * NUM_INPUTS]),
						.data_out(data_out[DATAW * (((SLICE_END - 1) >= SLICE_BEGIN ? SLICE_END - 1 : ((SLICE_END - 1) + ((SLICE_END - 1) >= SLICE_BEGIN ? ((SLICE_END - 1) - SLICE_BEGIN) + 1 : (SLICE_BEGIN - (SLICE_END - 1)) + 1)) - 1) - (((SLICE_END - 1) >= SLICE_BEGIN ? ((SLICE_END - 1) - SLICE_BEGIN) + 1 : (SLICE_BEGIN - (SLICE_END - 1)) + 1) - 1))+:DATAW * ((SLICE_END - 1) >= SLICE_BEGIN ? ((SLICE_END - 1) - SLICE_BEGIN) + 1 : (SLICE_BEGIN - (SLICE_END - 1)) + 1)]),
						.valid_out(valid_out[SLICE_END - 1:SLICE_BEGIN]),
						.ready_out(ready_out[SLICE_END - 1:SLICE_BEGIN]),
						.sel_out(sel_out_w[LOG_NUM_REQS2 * (s * NUM_INPUTS)+:LOG_NUM_REQS2 * NUM_INPUTS])
					);
				end
				genvar _gv_i_85;
				for (_gv_i_85 = 0; _gv_i_85 < NUM_INPUTS; _gv_i_85 = _gv_i_85 + 1) begin : g_sel_out
					localparam i = _gv_i_85;
					// Trace: src/VX_stream_arb.sv:214:17
					assign sel_out[i * NUM_REQS_W+:NUM_REQS_W] = {sel_tmp[i * LOG_NUM_REQS3+:LOG_NUM_REQS3], sel_out_w[((sel_tmp[i * LOG_NUM_REQS3+:LOG_NUM_REQS3] * NUM_INPUTS) + i) * LOG_NUM_REQS2+:LOG_NUM_REQS2]};
				end
			end
			else begin : g_arbiter
				// Trace: src/VX_stream_arb.sv:217:13
				wire [NUM_REQS - 1:0] arb_requests;
				// Trace: src/VX_stream_arb.sv:218:13
				wire arb_valid;
				// Trace: src/VX_stream_arb.sv:219:13
				wire [NUM_REQS_W - 1:0] arb_index;
				// Trace: src/VX_stream_arb.sv:220:13
				wire [NUM_REQS - 1:0] arb_onehot;
				// Trace: src/VX_stream_arb.sv:221:13
				wire arb_ready;
				genvar _gv_r_9;
				for (_gv_r_9 = 0; _gv_r_9 < NUM_REQS; _gv_r_9 = _gv_r_9 + 1) begin : g_requests
					localparam r = _gv_r_9;
					// Trace: src/VX_stream_arb.sv:223:17
					wire [NUM_INPUTS - 1:0] requests;
					genvar _gv_i_86;
					for (_gv_i_86 = 0; _gv_i_86 < NUM_INPUTS; _gv_i_86 = _gv_i_86 + 1) begin : g_i
						localparam i = _gv_i_86;
						// Trace: src/VX_stream_arb.sv:225:21
						localparam o = (r * NUM_INPUTS) + i;
						// Trace: src/VX_stream_arb.sv:226:21
						assign requests[i] = ready_out[o];
					end
					// Trace: src/VX_stream_arb.sv:228:17
					assign arb_requests[r] = |requests;
				end
				// Trace: src/VX_stream_arb.sv:230:13
				VX_generic_arbiter #(
					.NUM_REQS(NUM_REQS),
					.TYPE(ARBITER),
					.STICKY(STICKY)
				) arbiter(
					.clk(clk),
					.reset(reset),
					.requests(arb_requests),
					.grant_valid(arb_valid),
					.grant_index(arb_index),
					.grant_onehot(arb_onehot),
					.grant_ready(arb_ready)
				);
				// Trace: src/VX_stream_arb.sv:243:13
				wire [NUM_OUTPUTS - 1:0] valid_out_w;
				// Trace: src/VX_stream_arb.sv:244:13
				wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out_w;
				// Trace: src/VX_stream_arb.sv:245:13
				wire [NUM_OUTPUTS - 1:0] ready_out_w;
				genvar _gv_o_6;
				for (_gv_o_6 = 0; _gv_o_6 < NUM_OUTPUTS; _gv_o_6 = _gv_o_6 + 1) begin : g_data_out_w
					localparam o = _gv_o_6;
					// Trace: src/VX_stream_arb.sv:247:17
					localparam i = o % NUM_INPUTS;
					// Trace: src/VX_stream_arb.sv:248:17
					localparam r = o / NUM_INPUTS;
					// Trace: src/VX_stream_arb.sv:249:17
					assign valid_out_w[o] = valid_in[i] && arb_onehot[r];
					// Trace: src/VX_stream_arb.sv:250:17
					assign data_out_w[o * DATAW+:DATAW] = data_in[i * DATAW+:DATAW];
				end
				genvar _gv_i_87;
				for (_gv_i_87 = 0; _gv_i_87 < NUM_INPUTS; _gv_i_87 = _gv_i_87 + 1) begin : g_ready_in
					localparam i = _gv_i_87;
					// Trace: src/VX_stream_arb.sv:253:17
					wire [NUM_REQS - 1:0] ready_out_s;
					genvar _gv_r_10;
					for (_gv_r_10 = 0; _gv_r_10 < NUM_REQS; _gv_r_10 = _gv_r_10 + 1) begin : g_r
						localparam r = _gv_r_10;
						// Trace: src/VX_stream_arb.sv:255:21
						localparam o = (r * NUM_INPUTS) + i;
						// Trace: src/VX_stream_arb.sv:256:21
						assign ready_out_s[r] = ready_out_w[o];
					end
					// Trace: src/VX_stream_arb.sv:258:17
					assign ready_in[i] = (NUM_INPUTS == 1 ? arb_valid : |(ready_out_s & arb_onehot));
				end
				// Trace: src/VX_stream_arb.sv:260:13
				assign arb_ready = |valid_in;
				genvar _gv_o_7;
				for (_gv_o_7 = 0; _gv_o_7 < NUM_OUTPUTS; _gv_o_7 = _gv_o_7 + 1) begin : g_out_buf
					localparam o = _gv_o_7;
					// Trace: src/VX_stream_arb.sv:262:17
					VX_elastic_buffer #(
						.DATAW(DATAW),
						.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
						.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2)),
						.LUTRAM((OUT_BUF & 8) != 0)
					) out_buf(
						.clk(clk),
						.reset(reset),
						.valid_in(valid_out_w[o]),
						.ready_in(ready_out_w[o]),
						.data_in(data_out_w[o * DATAW+:DATAW]),
						.data_out(data_out[o * DATAW+:DATAW]),
						.valid_out(valid_out[o]),
						.ready_out(ready_out[o])
					);
				end
				genvar _gv_i_88;
				for (_gv_i_88 = 0; _gv_i_88 < NUM_INPUTS; _gv_i_88 = _gv_i_88 + 1) begin : g_sel_out
					localparam i = _gv_i_88;
					// Trace: src/VX_stream_arb.sv:279:17
					assign sel_out[i * NUM_REQS_W+:NUM_REQS_W] = arb_index;
				end
			end
		end
		else begin : g_passthru
			genvar _gv_o_8;
			for (_gv_o_8 = 0; _gv_o_8 < NUM_OUTPUTS; _gv_o_8 = _gv_o_8 + 1) begin : g_out_buf
				localparam o = _gv_o_8;
				// Trace: src/VX_stream_arb.sv:284:13
				VX_elastic_buffer #(
					.DATAW(DATAW),
					.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
					.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2)),
					.LUTRAM((OUT_BUF & 8) != 0)
				) out_buf(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_in[o]),
					.ready_in(ready_in[o]),
					.data_in(data_in[o * DATAW+:DATAW]),
					.data_out(data_out[o * DATAW+:DATAW]),
					.valid_out(valid_out[o]),
					.ready_out(ready_out[o])
				);
				// Trace: src/VX_stream_arb.sv:299:13
				assign sel_out[o * NUM_REQS_W+:NUM_REQS_W] = sv2v_cast_A9560_signed(0);
			end
		end
	endgenerate
endmodule
// removed interface: VX_dispatch_if
module VX_ipdom_stack (
	clk,
	reset,
	wid,
	d0,
	d1,
	rd_ptr,
	push,
	pop,
	q_val,
	q_idx,
	wr_ptr,
	empty,
	full
);
	// removed import VX_gpu_pkg::*;
	// Trace: src/VX_ipdom_stack.sv:2:15
	parameter WIDTH = 1;
	// Trace: src/VX_ipdom_stack.sv:3:15
	parameter DEPTH = 1;
	// Trace: src/VX_ipdom_stack.sv:4:15
	parameter ADDRW = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	// Trace: src/VX_ipdom_stack.sv:6:5
	input wire clk;
	// Trace: src/VX_ipdom_stack.sv:7:5
	input wire reset;
	// Trace: src/VX_ipdom_stack.sv:8:5
	localparam VX_gpu_pkg_NW_BITS = 2;
	localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
	input wire [1:0] wid;
	// Trace: src/VX_ipdom_stack.sv:9:5
	input wire [WIDTH - 1:0] d0;
	// Trace: src/VX_ipdom_stack.sv:10:5
	input wire [WIDTH - 1:0] d1;
	// Trace: src/VX_ipdom_stack.sv:11:5
	input wire [ADDRW - 1:0] rd_ptr;
	// Trace: src/VX_ipdom_stack.sv:12:5
	input wire push;
	// Trace: src/VX_ipdom_stack.sv:13:5
	input wire pop;
	// Trace: src/VX_ipdom_stack.sv:14:5
	output wire [WIDTH - 1:0] q_val;
	// Trace: src/VX_ipdom_stack.sv:15:5
	output wire q_idx;
	// Trace: src/VX_ipdom_stack.sv:16:5
	output wire [(4 * ADDRW) - 1:0] wr_ptr;
	// Trace: src/VX_ipdom_stack.sv:17:5
	output wire empty;
	// Trace: src/VX_ipdom_stack.sv:18:5
	output wire full;
	// Trace: src/VX_ipdom_stack.sv:20:5
	localparam BRAM_DATAW = 1 + (WIDTH * 2);
	// Trace: src/VX_ipdom_stack.sv:21:5
	localparam BRAM_SIZE = DEPTH * 4;
	// Trace: src/VX_ipdom_stack.sv:22:5
	localparam BRAW_ADDRW = (BRAM_SIZE > 1 ? $clog2(BRAM_SIZE) : 1);
	// Trace: src/VX_ipdom_stack.sv:23:5
	wire [(4 * ADDRW) - 1:0] wr_ptr_w;
	// Trace: src/VX_ipdom_stack.sv:24:5
	wire [3:0] empty_w;
	wire [3:0] full_w;
	// Trace: src/VX_ipdom_stack.sv:25:5
	genvar _gv_i_90;
	function automatic signed [ADDRW - 1:0] sv2v_cast_8BB5D_signed;
		input reg signed [ADDRW - 1:0] inp;
		sv2v_cast_8BB5D_signed = inp;
	endfunction
	function automatic [ADDRW - 1:0] sv2v_cast_8BB5D;
		input reg [ADDRW - 1:0] inp;
		sv2v_cast_8BB5D = inp;
	endfunction
	generate
		for (_gv_i_90 = 0; _gv_i_90 < 4; _gv_i_90 = _gv_i_90 + 1) begin : g_addressing
			localparam i = _gv_i_90;
			// Trace: src/VX_ipdom_stack.sv:26:9
			reg [ADDRW - 1:0] wr_ptr_r;
			// Trace: src/VX_ipdom_stack.sv:27:9
			reg empty_r;
			reg full_r;
			// Trace: src/VX_ipdom_stack.sv:28:9
			wire push_s = push && (wid == i);
			// Trace: src/VX_ipdom_stack.sv:29:9
			wire pop_s = pop && (wid == i);
			// Trace: src/VX_ipdom_stack.sv:33:9
			always @(posedge clk)
				// Trace: src/VX_ipdom_stack.sv:34:13
				if (reset) begin
					// Trace: src/VX_ipdom_stack.sv:35:17
					wr_ptr_r <= 1'sb0;
					// Trace: src/VX_ipdom_stack.sv:36:17
					empty_r <= 1;
					// Trace: src/VX_ipdom_stack.sv:37:17
					full_r <= 0;
				end
				else
					// Trace: src/VX_ipdom_stack.sv:39:17
					if (push_s) begin
						// Trace: src/VX_ipdom_stack.sv:40:21
						wr_ptr_r <= wr_ptr_r + sv2v_cast_8BB5D_signed(1);
						// Trace: src/VX_ipdom_stack.sv:41:21
						empty_r <= 0;
						// Trace: src/VX_ipdom_stack.sv:42:21
						full_r <= sv2v_cast_8BB5D_signed(DEPTH - 1) == wr_ptr_r;
					end
					else if (pop_s) begin
						// Trace: src/VX_ipdom_stack.sv:44:21
						wr_ptr_r <= wr_ptr_r - sv2v_cast_8BB5D(q_idx);
						// Trace: src/VX_ipdom_stack.sv:45:21
						empty_r <= (rd_ptr == 0) && q_idx;
						// Trace: src/VX_ipdom_stack.sv:46:21
						full_r <= 0;
					end
			// Trace: src/VX_ipdom_stack.sv:50:9
			assign wr_ptr_w[i * ADDRW+:ADDRW] = wr_ptr_r;
			// Trace: src/VX_ipdom_stack.sv:51:9
			assign empty_w[i] = empty_r;
			// Trace: src/VX_ipdom_stack.sv:52:9
			assign full_w[i] = full_r;
		end
	endgenerate
	// Trace: src/VX_ipdom_stack.sv:54:5
	wire [BRAW_ADDRW - 1:0] raddr;
	wire [BRAW_ADDRW - 1:0] waddr;
	// Trace: src/VX_ipdom_stack.sv:55:5
	generate
		if ((DEPTH > 1) && 1'd1) begin : g_DW
			// Trace: src/VX_ipdom_stack.sv:56:9
			assign waddr = (push ? {wr_ptr_w[wid * ADDRW+:ADDRW], wid} : {rd_ptr, wid});
			// Trace: src/VX_ipdom_stack.sv:57:9
			assign raddr = {rd_ptr, wid};
		end
		else if (DEPTH > 1) begin : g_D
			// Trace: src/VX_ipdom_stack.sv:59:9
			assign waddr = (push ? wr_ptr_w : rd_ptr);
			// Trace: src/VX_ipdom_stack.sv:60:9
			assign raddr = rd_ptr;
		end
		else begin : g_W
			// Trace: src/VX_ipdom_stack.sv:62:9
			assign waddr = (push ? wid : wid);
			// Trace: src/VX_ipdom_stack.sv:63:9
			assign raddr = 0;
		end
	endgenerate
	// Trace: src/VX_ipdom_stack.sv:68:5
	wire [WIDTH - 1:0] q0;
	wire [WIDTH - 1:0] q1;
	// Trace: src/VX_ipdom_stack.sv:69:5
	VX_dp_ram #(
		.DATAW(BRAM_DATAW),
		.SIZE(BRAM_SIZE),
		.RDW_MODE("R"),
		.RADDR_REG(1)
	) ipdom_store(
		.clk(clk),
		.reset(reset),
		.read(pop),
		.write(push || pop),
		.wren(1'b1),
		.waddr(waddr),
		.raddr(raddr),
		.wdata((push ? {1'b0, d1, d0} : {1'b1, q1, q0})),
		.rdata({q_idx, q1, q0})
	);
	// Trace: src/VX_ipdom_stack.sv:85:5
	assign q_val = (q_idx ? q0 : q1);
	// Trace: src/VX_ipdom_stack.sv:86:5
	assign wr_ptr = wr_ptr_w;
	// Trace: src/VX_ipdom_stack.sv:87:5
	assign empty = empty_w[wid];
	// Trace: src/VX_ipdom_stack.sv:88:5
	assign full = full_w[wid];
endmodule
// removed module with interface ports: VX_dispatch
module Vortex (
	clk,
	reset,
	mem_req_valid,
	mem_req_rw,
	mem_req_byteen,
	mem_req_addr,
	mem_req_data,
	mem_req_tag,
	mem_req_ready,
	mem_rsp_valid,
	mem_rsp_data,
	mem_rsp_tag,
	mem_rsp_ready,
	dcr_wr_valid,
	dcr_wr_addr,
	dcr_wr_data,
	busy
);
	// removed import VX_gpu_pkg::*;
	// Trace: src/Vortex.sv:2:5
	input wire clk;
	// Trace: src/Vortex.sv:3:5
	input wire reset;
	// Trace: src/Vortex.sv:4:5
	localparam VX_gpu_pkg_DCACHE_WORD_SIZE = 16;
	localparam VX_gpu_pkg_XLENB = 4;
	localparam VX_gpu_pkg_LSU_WORD_SIZE = VX_gpu_pkg_XLENB;
	localparam VX_gpu_pkg_DCACHE_CHANNELS = 1;
	localparam VX_gpu_pkg_DCACHE_NUM_REQS = 1;
	localparam VX_gpu_pkg_NUM_SOCKETS = 1;
	localparam VX_gpu_pkg_L2_NUM_REQS = 1;
	localparam VX_gpu_pkg_L3_NUM_REQS = 1;
	localparam VX_gpu_pkg_VX_MEM_PORTS = VX_gpu_pkg_L3_NUM_REQS;
	output wire [0:0] mem_req_valid;
	// Trace: src/Vortex.sv:5:5
	output wire [0:0] mem_req_rw;
	// Trace: src/Vortex.sv:6:5
	localparam VX_gpu_pkg_VX_MEM_BYTEEN_WIDTH = 64;
	output wire [63:0] mem_req_byteen;
	// Trace: src/Vortex.sv:7:5
	localparam VX_gpu_pkg_VX_MEM_ADDR_WIDTH = 26;
	output wire [25:0] mem_req_addr;
	// Trace: src/Vortex.sv:8:5
	localparam VX_gpu_pkg_VX_MEM_DATA_WIDTH = 512;
	output wire [511:0] mem_req_data;
	// Trace: src/Vortex.sv:9:5
	localparam VX_gpu_pkg_DCACHE_LINE_SIZE = 64;
	localparam VX_gpu_pkg_DCACHE_MERGED_REQS = 1;
	localparam VX_gpu_pkg_DCACHE_MEM_BATCHES = 1;
	localparam VX_gpu_pkg_DCACHE_TAG_ID_BITS = 2;
	localparam VX_gpu_pkg_UUID_WIDTH = 1;
	localparam VX_gpu_pkg_DCACHE_TAG_WIDTH = 3;
	localparam VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH = 6;
	localparam VX_gpu_pkg_ICACHE_MEM_TAG_WIDTH = 5;
	localparam VX_gpu_pkg_L1_MEM_TAG_WIDTH = VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH;
	localparam VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH = 7;
	localparam VX_gpu_pkg_L2_TAG_WIDTH = VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH;
	localparam VX_gpu_pkg_L2_WORD_SIZE = 64;
	localparam VX_gpu_pkg_L2_MEM_TAG_WIDTH = 7;
	localparam VX_gpu_pkg_L3_TAG_WIDTH = VX_gpu_pkg_L2_MEM_TAG_WIDTH;
	localparam VX_gpu_pkg_L3_WORD_SIZE = 64;
	localparam VX_gpu_pkg_L3_MEM_TAG_WIDTH = 7;
	localparam VX_gpu_pkg_VX_MEM_TAG_WIDTH = VX_gpu_pkg_L3_MEM_TAG_WIDTH;
	output wire [6:0] mem_req_tag;
	// Trace: src/Vortex.sv:10:5
	input wire [0:0] mem_req_ready;
	// Trace: src/Vortex.sv:11:5
	input wire [0:0] mem_rsp_valid;
	// Trace: src/Vortex.sv:12:5
	input wire [511:0] mem_rsp_data;
	// Trace: src/Vortex.sv:13:5
	input wire [6:0] mem_rsp_tag;
	// Trace: src/Vortex.sv:14:5
	output wire [0:0] mem_rsp_ready;
	// Trace: src/Vortex.sv:15:5
	input wire dcr_wr_valid;
	// Trace: src/Vortex.sv:16:5
	localparam VX_gpu_pkg_VX_DCR_ADDR_WIDTH = 12;
	input wire [11:0] dcr_wr_addr;
	// Trace: src/Vortex.sv:17:5
	localparam VX_gpu_pkg_VX_DCR_DATA_WIDTH = 32;
	input wire [31:0] dcr_wr_data;
	// Trace: src/Vortex.sv:18:5
	output wire busy;
	// Trace: src/Vortex.sv:20:5
	// expanded interface instance: per_cluster_mem_bus_if
	localparam _param_CA4E3_DATA_SIZE = 64;
	localparam _param_CA4E3_TAG_WIDTH = VX_gpu_pkg_L2_MEM_TAG_WIDTH;
	genvar _arr_CA4E3;
	generate
		for (_arr_CA4E3 = 0; _arr_CA4E3 <= 0; _arr_CA4E3 = _arr_CA4E3 + 1) begin : per_cluster_mem_bus_if
			// removed import VX_gpu_pkg::*;
			// Trace: src/VX_mem_bus_if.sv:2:15
			localparam DATA_SIZE = _param_CA4E3_DATA_SIZE;
			// Trace: src/VX_mem_bus_if.sv:3:15
			localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
			localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
			localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
			// Trace: src/VX_mem_bus_if.sv:4:15
			localparam TAG_WIDTH = _param_CA4E3_TAG_WIDTH;
			// Trace: src/VX_mem_bus_if.sv:5:15
			localparam MEM_ADDR_WIDTH = 32;
			// Trace: src/VX_mem_bus_if.sv:6:15
			localparam ADDR_WIDTH = 26;
			// Trace: src/VX_mem_bus_if.sv:8:5
			localparam VX_gpu_pkg_UUID_WIDTH = 1;
			// removed localparam type tag_t
			// Trace: src/VX_mem_bus_if.sv:12:5
			// removed localparam type req_data_t
			// Trace: src/VX_mem_bus_if.sv:20:5
			// removed localparam type rsp_data_t
			// Trace: src/VX_mem_bus_if.sv:24:5
			wire req_valid;
			// Trace: src/VX_mem_bus_if.sv:25:5
			wire [612:0] req_data;
			// Trace: src/VX_mem_bus_if.sv:26:5
			wire req_ready;
			// Trace: src/VX_mem_bus_if.sv:27:5
			wire rsp_valid;
			// Trace: src/VX_mem_bus_if.sv:28:5
			wire [518:0] rsp_data;
			// Trace: src/VX_mem_bus_if.sv:29:5
			wire rsp_ready;
			// Trace: src/VX_mem_bus_if.sv:30:5
			// Trace: src/VX_mem_bus_if.sv:38:5
		end
	endgenerate
	// Trace: src/Vortex.sv:24:5
	// expanded interface instance: mem_bus_if
	localparam _param_4F26C_DATA_SIZE = 64;
	localparam _param_4F26C_TAG_WIDTH = VX_gpu_pkg_L3_MEM_TAG_WIDTH;
	genvar _arr_4F26C;
	generate
		for (_arr_4F26C = 0; _arr_4F26C <= 0; _arr_4F26C = _arr_4F26C + 1) begin : mem_bus_if
			// removed import VX_gpu_pkg::*;
			// Trace: src/VX_mem_bus_if.sv:2:15
			localparam DATA_SIZE = _param_4F26C_DATA_SIZE;
			// Trace: src/VX_mem_bus_if.sv:3:15
			localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
			localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
			localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
			// Trace: src/VX_mem_bus_if.sv:4:15
			localparam TAG_WIDTH = _param_4F26C_TAG_WIDTH;
			// Trace: src/VX_mem_bus_if.sv:5:15
			localparam MEM_ADDR_WIDTH = 32;
			// Trace: src/VX_mem_bus_if.sv:6:15
			localparam ADDR_WIDTH = 26;
			// Trace: src/VX_mem_bus_if.sv:8:5
			localparam VX_gpu_pkg_UUID_WIDTH = 1;
			// removed localparam type tag_t
			// Trace: src/VX_mem_bus_if.sv:12:5
			// removed localparam type req_data_t
			// Trace: src/VX_mem_bus_if.sv:20:5
			// removed localparam type rsp_data_t
			// Trace: src/VX_mem_bus_if.sv:24:5
			wire req_valid;
			// Trace: src/VX_mem_bus_if.sv:25:5
			wire [612:0] req_data;
			// Trace: src/VX_mem_bus_if.sv:26:5
			wire req_ready;
			// Trace: src/VX_mem_bus_if.sv:27:5
			wire rsp_valid;
			// Trace: src/VX_mem_bus_if.sv:28:5
			wire [518:0] rsp_data;
			// Trace: src/VX_mem_bus_if.sv:29:5
			wire rsp_ready;
			// Trace: src/VX_mem_bus_if.sv:30:5
			// Trace: src/VX_mem_bus_if.sv:38:5
		end
	endgenerate
	// Trace: src/Vortex.sv:28:5
	wire [0:0] l3_reset;
	// Trace: src/Vortex.sv:29:5
	VX_reset_relay #(
		.N(1),
		.MAX_FANOUT(0)
	) __l3_reset(
		.clk(clk),
		.reset(reset),
		.reset_o(l3_reset)
	);
	// Trace: src/Vortex.sv:34:5
	// expanded module instance: l3cache
	localparam _bbase_56375_core_bus_if = 0;
	localparam _bbase_56375_mem_bus_if = 0;
	localparam _param_56375_INSTANCE_ID = "l3cache";
	localparam _param_56375_CACHE_SIZE = 2097152;
	localparam _param_56375_LINE_SIZE = 64;
	localparam _param_56375_NUM_BANKS = VX_gpu_pkg_L3_NUM_REQS;
	localparam _param_56375_NUM_WAYS = 8;
	localparam _param_56375_WORD_SIZE = VX_gpu_pkg_L3_WORD_SIZE;
	localparam _param_56375_NUM_REQS = VX_gpu_pkg_L3_NUM_REQS;
	localparam _param_56375_MEM_PORTS = VX_gpu_pkg_L3_NUM_REQS;
	localparam _param_56375_CRSQ_SIZE = 2;
	localparam _param_56375_MSHR_SIZE = 16;
	localparam _param_56375_MRSQ_SIZE = 4;
	localparam _param_56375_MREQ_SIZE = 4;
	localparam _param_56375_TAG_WIDTH = VX_gpu_pkg_L2_MEM_TAG_WIDTH;
	localparam _param_56375_WRITE_ENABLE = 1;
	localparam _param_56375_WRITEBACK = 0;
	localparam _param_56375_DIRTY_BYTES = 0;
	localparam _param_56375_REPL_POLICY = 1;
	localparam _param_56375_CORE_OUT_BUF = 3;
	localparam _param_56375_MEM_OUT_BUF = 3;
	localparam _param_56375_NC_ENABLE = 1;
	localparam _param_56375_PASSTHRU = 1'd1;
	function automatic [6:0] sv2v_cast_7;
		input reg [6:0] inp;
		sv2v_cast_7 = inp;
	endfunction
	generate
		if (1) begin : l3cache
			// removed import VX_gpu_pkg::*;
			// Trace: src/VX_cache_wrap.sv:2:15
			localparam INSTANCE_ID = _param_56375_INSTANCE_ID;
			// Trace: src/VX_cache_wrap.sv:3:15
			localparam TAG_SEL_IDX = 0;
			// Trace: src/VX_cache_wrap.sv:4:15
			localparam NUM_REQS = _param_56375_NUM_REQS;
			// Trace: src/VX_cache_wrap.sv:5:15
			localparam MEM_PORTS = _param_56375_MEM_PORTS;
			// Trace: src/VX_cache_wrap.sv:6:15
			localparam CACHE_SIZE = _param_56375_CACHE_SIZE;
			// Trace: src/VX_cache_wrap.sv:7:15
			localparam LINE_SIZE = _param_56375_LINE_SIZE;
			// Trace: src/VX_cache_wrap.sv:8:15
			localparam NUM_BANKS = _param_56375_NUM_BANKS;
			// Trace: src/VX_cache_wrap.sv:9:15
			localparam NUM_WAYS = _param_56375_NUM_WAYS;
			// Trace: src/VX_cache_wrap.sv:10:15
			localparam WORD_SIZE = _param_56375_WORD_SIZE;
			// Trace: src/VX_cache_wrap.sv:11:15
			localparam CRSQ_SIZE = _param_56375_CRSQ_SIZE;
			// Trace: src/VX_cache_wrap.sv:12:15
			localparam MSHR_SIZE = _param_56375_MSHR_SIZE;
			// Trace: src/VX_cache_wrap.sv:13:15
			localparam MRSQ_SIZE = _param_56375_MRSQ_SIZE;
			// Trace: src/VX_cache_wrap.sv:14:15
			localparam MREQ_SIZE = _param_56375_MREQ_SIZE;
			// Trace: src/VX_cache_wrap.sv:15:15
			localparam WRITE_ENABLE = _param_56375_WRITE_ENABLE;
			// Trace: src/VX_cache_wrap.sv:16:15
			localparam WRITEBACK = _param_56375_WRITEBACK;
			// Trace: src/VX_cache_wrap.sv:17:15
			localparam DIRTY_BYTES = _param_56375_DIRTY_BYTES;
			// Trace: src/VX_cache_wrap.sv:18:15
			localparam REPL_POLICY = _param_56375_REPL_POLICY;
			// Trace: src/VX_cache_wrap.sv:19:15
			localparam VX_gpu_pkg_UUID_WIDTH = 1;
			localparam TAG_WIDTH = _param_56375_TAG_WIDTH;
			// Trace: src/VX_cache_wrap.sv:20:15
			localparam NC_ENABLE = _param_56375_NC_ENABLE;
			// Trace: src/VX_cache_wrap.sv:21:15
			localparam PASSTHRU = _param_56375_PASSTHRU;
			// Trace: src/VX_cache_wrap.sv:22:15
			localparam CORE_OUT_BUF = _param_56375_CORE_OUT_BUF;
			// Trace: src/VX_cache_wrap.sv:23:15
			localparam MEM_OUT_BUF = _param_56375_MEM_OUT_BUF;
			// Trace: src/VX_cache_wrap.sv:25:5
			wire clk;
			// Trace: src/VX_cache_wrap.sv:26:5
			wire reset;
			// Trace: src/VX_cache_wrap.sv:27:5
			localparam _mbase_core_bus_if = 0;
			// Trace: src/VX_cache_wrap.sv:28:5
			localparam _mbase_mem_bus_if = 0;
			// Trace: src/VX_cache_wrap.sv:30:5
			localparam CACHE_MEM_TAG_WIDTH = 5;
			// Trace: src/VX_cache_wrap.sv:32:5
			localparam BYPASS_TAG_WIDTH = 7;
			// Trace: src/VX_cache_wrap.sv:34:5
			localparam NC_TAG_WIDTH = 8;
			// Trace: src/VX_cache_wrap.sv:35:5
			localparam MEM_TAG_WIDTH = (PASSTHRU ? BYPASS_TAG_WIDTH : (NC_ENABLE ? NC_TAG_WIDTH : CACHE_MEM_TAG_WIDTH));
			// Trace: src/VX_cache_wrap.sv:36:5
			localparam BYPASS_ENABLE = 1'd1;
			// Trace: src/VX_cache_wrap.sv:37:5
			// expanded interface instance: core_bus_cache_if
			localparam _param_24C1C_DATA_SIZE = WORD_SIZE;
			localparam _param_24C1C_TAG_WIDTH = TAG_WIDTH;
			genvar _arr_24C1C;
			for (_arr_24C1C = 0; _arr_24C1C <= 0; _arr_24C1C = _arr_24C1C + 1) begin : core_bus_cache_if
				// removed import VX_gpu_pkg::*;
				// Trace: src/VX_mem_bus_if.sv:2:15
				localparam DATA_SIZE = _param_24C1C_DATA_SIZE;
				// Trace: src/VX_mem_bus_if.sv:3:15
				localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
				localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
				localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
				// Trace: src/VX_mem_bus_if.sv:4:15
				localparam TAG_WIDTH = _param_24C1C_TAG_WIDTH;
				// Trace: src/VX_mem_bus_if.sv:5:15
				localparam MEM_ADDR_WIDTH = 32;
				// Trace: src/VX_mem_bus_if.sv:6:15
				localparam ADDR_WIDTH = 26;
				// Trace: src/VX_mem_bus_if.sv:8:5
				localparam VX_gpu_pkg_UUID_WIDTH = 1;
				// removed localparam type tag_t
				// Trace: src/VX_mem_bus_if.sv:12:5
				// removed localparam type req_data_t
				// Trace: src/VX_mem_bus_if.sv:20:5
				// removed localparam type rsp_data_t
				// Trace: src/VX_mem_bus_if.sv:24:5
				wire req_valid;
				// Trace: src/VX_mem_bus_if.sv:25:5
				wire [612:0] req_data;
				// Trace: src/VX_mem_bus_if.sv:26:5
				wire req_ready;
				// Trace: src/VX_mem_bus_if.sv:27:5
				wire rsp_valid;
				// Trace: src/VX_mem_bus_if.sv:28:5
				wire [518:0] rsp_data;
				// Trace: src/VX_mem_bus_if.sv:29:5
				wire rsp_ready;
				// Trace: src/VX_mem_bus_if.sv:30:5
				// Trace: src/VX_mem_bus_if.sv:38:5
			end
			// Trace: src/VX_cache_wrap.sv:41:5
			// expanded interface instance: mem_bus_cache_if
			localparam _param_D895D_DATA_SIZE = LINE_SIZE;
			localparam _param_D895D_TAG_WIDTH = CACHE_MEM_TAG_WIDTH;
			genvar _arr_D895D;
			for (_arr_D895D = 0; _arr_D895D <= 0; _arr_D895D = _arr_D895D + 1) begin : mem_bus_cache_if
				// removed import VX_gpu_pkg::*;
				// Trace: src/VX_mem_bus_if.sv:2:15
				localparam DATA_SIZE = _param_D895D_DATA_SIZE;
				// Trace: src/VX_mem_bus_if.sv:3:15
				localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
				localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
				localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
				// Trace: src/VX_mem_bus_if.sv:4:15
				localparam TAG_WIDTH = _param_D895D_TAG_WIDTH;
				// Trace: src/VX_mem_bus_if.sv:5:15
				localparam MEM_ADDR_WIDTH = 32;
				// Trace: src/VX_mem_bus_if.sv:6:15
				localparam ADDR_WIDTH = 26;
				// Trace: src/VX_mem_bus_if.sv:8:5
				localparam VX_gpu_pkg_UUID_WIDTH = 1;
				// removed localparam type tag_t
				// Trace: src/VX_mem_bus_if.sv:12:5
				// removed localparam type req_data_t
				// Trace: src/VX_mem_bus_if.sv:20:5
				// removed localparam type rsp_data_t
				// Trace: src/VX_mem_bus_if.sv:24:5
				wire req_valid;
				// Trace: src/VX_mem_bus_if.sv:25:5
				wire [610:0] req_data;
				// Trace: src/VX_mem_bus_if.sv:26:5
				wire req_ready;
				// Trace: src/VX_mem_bus_if.sv:27:5
				wire rsp_valid;
				// Trace: src/VX_mem_bus_if.sv:28:5
				wire [516:0] rsp_data;
				// Trace: src/VX_mem_bus_if.sv:29:5
				wire rsp_ready;
				// Trace: src/VX_mem_bus_if.sv:30:5
				// Trace: src/VX_mem_bus_if.sv:38:5
			end
			// Trace: src/VX_cache_wrap.sv:45:5
			// expanded interface instance: mem_bus_tmp_if
			localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
			localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH;
			genvar _arr_4FE36;
			for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
				// removed import VX_gpu_pkg::*;
				// Trace: src/VX_mem_bus_if.sv:2:15
				localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
				// Trace: src/VX_mem_bus_if.sv:3:15
				localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
				localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
				localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
				// Trace: src/VX_mem_bus_if.sv:4:15
				localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
				// Trace: src/VX_mem_bus_if.sv:5:15
				localparam MEM_ADDR_WIDTH = 32;
				// Trace: src/VX_mem_bus_if.sv:6:15
				localparam ADDR_WIDTH = 26;
				// Trace: src/VX_mem_bus_if.sv:8:5
				localparam VX_gpu_pkg_UUID_WIDTH = 1;
				// removed localparam type tag_t
				// Trace: src/VX_mem_bus_if.sv:12:5
				// removed localparam type req_data_t
				// Trace: src/VX_mem_bus_if.sv:20:5
				// removed localparam type rsp_data_t
				// Trace: src/VX_mem_bus_if.sv:24:5
				wire req_valid;
				// Trace: src/VX_mem_bus_if.sv:25:5
				wire [(606 + (_param_4FE36_TAG_WIDTH + 0)) - 1:0] req_data;
				// Trace: src/VX_mem_bus_if.sv:26:5
				wire req_ready;
				// Trace: src/VX_mem_bus_if.sv:27:5
				wire rsp_valid;
				// Trace: src/VX_mem_bus_if.sv:28:5
				wire [(512 + (_param_4FE36_TAG_WIDTH + 0)) - 1:0] rsp_data;
				// Trace: src/VX_mem_bus_if.sv:29:5
				wire rsp_ready;
				// Trace: src/VX_mem_bus_if.sv:30:5
				// Trace: src/VX_mem_bus_if.sv:38:5
			end
			// Trace: src/VX_cache_wrap.sv:49:5
			if (BYPASS_ENABLE) begin : g_bypass
				// Trace: src/VX_cache_wrap.sv:50:9
				// expanded module instance: cache_bypass
				localparam _bbase_714AA_core_bus_in_if = 0;
				localparam _bbase_714AA_core_bus_out_if = 0;
				localparam _bbase_714AA_mem_bus_in_if = 0;
				localparam _bbase_714AA_mem_bus_out_if = 0;
				localparam _param_714AA_NUM_REQS = NUM_REQS;
				localparam _param_714AA_MEM_PORTS = MEM_PORTS;
				localparam _param_714AA_TAG_SEL_IDX = TAG_SEL_IDX;
				localparam _param_714AA_CACHE_ENABLE = !PASSTHRU;
				localparam _param_714AA_WORD_SIZE = WORD_SIZE;
				localparam _param_714AA_LINE_SIZE = LINE_SIZE;
				localparam _param_714AA_CORE_ADDR_WIDTH = 26;
				localparam _param_714AA_CORE_TAG_WIDTH = TAG_WIDTH;
				localparam _param_714AA_MEM_ADDR_WIDTH = 26;
				localparam _param_714AA_MEM_TAG_IN_WIDTH = CACHE_MEM_TAG_WIDTH;
				localparam _param_714AA_CORE_OUT_BUF = CORE_OUT_BUF;
				localparam _param_714AA_MEM_OUT_BUF = MEM_OUT_BUF;
				if (1) begin : cache_bypass
					// removed import VX_gpu_pkg::*;
					// Trace: src/VX_cache_bypass.sv:2:15
					localparam NUM_REQS = _param_714AA_NUM_REQS;
					// Trace: src/VX_cache_bypass.sv:3:15
					localparam MEM_PORTS = _param_714AA_MEM_PORTS;
					// Trace: src/VX_cache_bypass.sv:4:15
					localparam TAG_SEL_IDX = _param_714AA_TAG_SEL_IDX;
					// Trace: src/VX_cache_bypass.sv:5:15
					localparam CACHE_ENABLE = _param_714AA_CACHE_ENABLE;
					// Trace: src/VX_cache_bypass.sv:6:15
					localparam WORD_SIZE = _param_714AA_WORD_SIZE;
					// Trace: src/VX_cache_bypass.sv:7:15
					localparam LINE_SIZE = _param_714AA_LINE_SIZE;
					// Trace: src/VX_cache_bypass.sv:8:15
					localparam CORE_ADDR_WIDTH = _param_714AA_CORE_ADDR_WIDTH;
					// Trace: src/VX_cache_bypass.sv:9:15
					localparam CORE_TAG_WIDTH = _param_714AA_CORE_TAG_WIDTH;
					// Trace: src/VX_cache_bypass.sv:10:15
					localparam MEM_ADDR_WIDTH = _param_714AA_MEM_ADDR_WIDTH;
					// Trace: src/VX_cache_bypass.sv:11:15
					localparam MEM_TAG_IN_WIDTH = _param_714AA_MEM_TAG_IN_WIDTH;
					// Trace: src/VX_cache_bypass.sv:12:15
					localparam CORE_OUT_BUF = _param_714AA_CORE_OUT_BUF;
					// Trace: src/VX_cache_bypass.sv:13:15
					localparam MEM_OUT_BUF = _param_714AA_MEM_OUT_BUF;
					// Trace: src/VX_cache_bypass.sv:15:5
					wire clk;
					// Trace: src/VX_cache_bypass.sv:16:5
					wire reset;
					// Trace: src/VX_cache_bypass.sv:17:5
					localparam _mbase_core_bus_in_if = 0;
					// Trace: src/VX_cache_bypass.sv:18:5
					localparam _mbase_core_bus_out_if = 0;
					// Trace: src/VX_cache_bypass.sv:19:5
					localparam _mbase_mem_bus_in_if = 0;
					// Trace: src/VX_cache_bypass.sv:20:5
					localparam _mbase_mem_bus_out_if = 0;
					// Trace: src/VX_cache_bypass.sv:22:5
					localparam DIRECT_PASSTHRU = (!CACHE_ENABLE && 1'd1) && 1'd1;
					// Trace: src/VX_cache_bypass.sv:23:5
					localparam CORE_DATA_WIDTH = 512;
					// Trace: src/VX_cache_bypass.sv:24:5
					localparam WORDS_PER_LINE = 1;
					// Trace: src/VX_cache_bypass.sv:25:5
					localparam WSEL_BITS = 0;
					// Trace: src/VX_cache_bypass.sv:26:5
					localparam VX_gpu_pkg_UUID_WIDTH = 1;
					localparam CORE_TAG_ID_WIDTH = 6;
					// Trace: src/VX_cache_bypass.sv:27:5
					localparam MEM_TAG_ID_WIDTH = 6;
					// Trace: src/VX_cache_bypass.sv:28:5
					localparam MEM_TAG_NC1_WIDTH = 7;
					// Trace: src/VX_cache_bypass.sv:29:5
					localparam MEM_TAG_NC2_WIDTH = 7;
					// Trace: src/VX_cache_bypass.sv:30:5
					localparam MEM_TAG_OUT_WIDTH = (CACHE_ENABLE ? MEM_TAG_NC2_WIDTH : MEM_TAG_NC2_WIDTH);
					// Trace: src/VX_cache_bypass.sv:31:5
					// expanded interface instance: core_bus_nc_switch_if
					localparam _param_95306_DATA_SIZE = WORD_SIZE;
					localparam _param_95306_TAG_WIDTH = CORE_TAG_WIDTH;
					genvar _arr_95306;
					for (_arr_95306 = 0; _arr_95306 <= (((CACHE_ENABLE ? 2 : 1) * NUM_REQS) - 1); _arr_95306 = _arr_95306 + 1) begin : core_bus_nc_switch_if
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_95306_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
						localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
						localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_95306_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:8:5
						localparam VX_gpu_pkg_UUID_WIDTH = 1;
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:12:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:20:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:24:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire [612:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire [518:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:30:5
						// Trace: src/VX_mem_bus_if.sv:38:5
					end
					// Trace: src/VX_cache_bypass.sv:35:5
					wire [0:0] core_req_nc_sel;
					// Trace: src/VX_cache_bypass.sv:36:5
					genvar _gv_i_56;
					localparam VX_gpu_pkg_MEM_REQ_FLAG_IO = 1;
					for (_gv_i_56 = 0; _gv_i_56 < NUM_REQS; _gv_i_56 = _gv_i_56 + 1) begin : g_core_req_is_nc
						localparam i = _gv_i_56;
						if (CACHE_ENABLE) begin : g_cache
							// Trace: src/VX_cache_bypass.sv:38:13
							assign core_req_nc_sel[i] = ~Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_in_if].req_data[8];
						end
						else begin : g_no_cache
							// Trace: src/VX_cache_bypass.sv:40:13
							assign core_req_nc_sel[i] = 1'b0;
						end
					end
					// Trace: src/VX_cache_bypass.sv:43:5
					// expanded module instance: core_bus_nc_switch
					localparam _bbase_69FDB_bus_in_if = 0;
					localparam _bbase_69FDB_bus_out_if = 0;
					localparam _param_69FDB_NUM_INPUTS = NUM_REQS;
					localparam _param_69FDB_NUM_OUTPUTS = (CACHE_ENABLE ? 2 : 1) * NUM_REQS;
					localparam _param_69FDB_DATA_SIZE = WORD_SIZE;
					localparam _param_69FDB_TAG_WIDTH = CORE_TAG_WIDTH;
					localparam _param_69FDB_ARBITER = "R";
					localparam _param_69FDB_REQ_OUT_BUF = 0;
					localparam _param_69FDB_RSP_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
					if (1) begin : core_bus_nc_switch
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_mem_switch.sv:2:15
						localparam NUM_INPUTS = _param_69FDB_NUM_INPUTS;
						// Trace: src/VX_mem_switch.sv:3:15
						localparam NUM_OUTPUTS = _param_69FDB_NUM_OUTPUTS;
						// Trace: src/VX_mem_switch.sv:4:15
						localparam DATA_SIZE = _param_69FDB_DATA_SIZE;
						// Trace: src/VX_mem_switch.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_switch.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_switch.sv:7:15
						localparam TAG_WIDTH = _param_69FDB_TAG_WIDTH;
						// Trace: src/VX_mem_switch.sv:8:15
						localparam REQ_OUT_BUF = _param_69FDB_REQ_OUT_BUF;
						// Trace: src/VX_mem_switch.sv:9:15
						localparam RSP_OUT_BUF = _param_69FDB_RSP_OUT_BUF;
						// Trace: src/VX_mem_switch.sv:10:15
						localparam ARBITER = _param_69FDB_ARBITER;
						// Trace: src/VX_mem_switch.sv:11:15
						localparam NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? ((NUM_INPUTS + NUM_OUTPUTS) - 1) / NUM_OUTPUTS : ((NUM_OUTPUTS + NUM_INPUTS) - 1) / NUM_INPUTS);
						// Trace: src/VX_mem_switch.sv:12:15
						localparam SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
						// Trace: src/VX_mem_switch.sv:13:15
						localparam LOG_NUM_REQS = $clog2(NUM_REQS);
						// Trace: src/VX_mem_switch.sv:15:5
						wire clk;
						// Trace: src/VX_mem_switch.sv:16:5
						wire reset;
						// Trace: src/VX_mem_switch.sv:17:5
						wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] bus_sel;
						// Trace: src/VX_mem_switch.sv:18:5
						localparam _mbase_bus_in_if = 0;
						// Trace: src/VX_mem_switch.sv:19:5
						localparam _mbase_bus_out_if = 0;
						// Trace: src/VX_mem_switch.sv:21:5
						localparam DATA_WIDTH = 512;
						// Trace: src/VX_mem_switch.sv:22:5
						localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
						localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
						localparam REQ_DATAW = 613;
						// Trace: src/VX_mem_switch.sv:23:5
						localparam RSP_DATAW = 519;
						// Trace: src/VX_mem_switch.sv:24:5
						wire [0:0] req_valid_in;
						// Trace: src/VX_mem_switch.sv:25:5
						wire [612:0] req_data_in;
						// Trace: src/VX_mem_switch.sv:26:5
						wire [0:0] req_ready_in;
						// Trace: src/VX_mem_switch.sv:27:5
						wire [NUM_OUTPUTS - 1:0] req_valid_out;
						// Trace: src/VX_mem_switch.sv:28:5
						wire [(NUM_OUTPUTS * 613) - 1:0] req_data_out;
						// Trace: src/VX_mem_switch.sv:29:5
						wire [NUM_OUTPUTS - 1:0] req_ready_out;
						// Trace: src/VX_mem_switch.sv:30:5
						genvar _gv_i_109;
						for (_gv_i_109 = 0; _gv_i_109 < NUM_INPUTS; _gv_i_109 = _gv_i_109 + 1) begin : g_req_data_in
							localparam i = _gv_i_109;
							// Trace: src/VX_mem_switch.sv:31:9
							assign req_valid_in[i] = Vortex.per_cluster_mem_bus_if[i + _mbase_bus_in_if].req_valid;
							// Trace: src/VX_mem_switch.sv:32:9
							assign req_data_in[i * 613+:613] = Vortex.per_cluster_mem_bus_if[i + _mbase_bus_in_if].req_data;
							// Trace: src/VX_mem_switch.sv:33:9
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
						end
						// Trace: src/VX_mem_switch.sv:35:5
						VX_stream_switch #(
							.NUM_INPUTS(NUM_INPUTS),
							.NUM_OUTPUTS(NUM_OUTPUTS),
							.DATAW(REQ_DATAW),
							.OUT_BUF(REQ_OUT_BUF)
						) req_switch(
							.clk(clk),
							.reset(reset),
							.sel_in(bus_sel),
							.valid_in(req_valid_in),
							.data_in(req_data_in),
							.ready_in(req_ready_in),
							.valid_out(req_valid_out),
							.data_out(req_data_out),
							.ready_out(req_ready_out)
						);
						// Trace: src/VX_mem_switch.sv:51:5
						genvar _gv_i_110;
						for (_gv_i_110 = 0; _gv_i_110 < NUM_OUTPUTS; _gv_i_110 = _gv_i_110 + 1) begin : g_req_data_out
							localparam i = _gv_i_110;
							// Trace: src/VX_mem_switch.sv:52:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
							// Trace: src/VX_mem_switch.sv:53:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_data = req_data_out[i * 613+:613];
							// Trace: src/VX_mem_switch.sv:54:9
							assign req_ready_out[i] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_ready;
						end
						// Trace: src/VX_mem_switch.sv:56:5
						wire [NUM_OUTPUTS - 1:0] rsp_valid_in;
						// Trace: src/VX_mem_switch.sv:57:5
						wire [(NUM_OUTPUTS * 519) - 1:0] rsp_data_in;
						// Trace: src/VX_mem_switch.sv:58:5
						wire [NUM_OUTPUTS - 1:0] rsp_ready_in;
						// Trace: src/VX_mem_switch.sv:59:5
						wire [0:0] rsp_valid_out;
						// Trace: src/VX_mem_switch.sv:60:5
						wire [518:0] rsp_data_out;
						// Trace: src/VX_mem_switch.sv:61:5
						wire [0:0] rsp_ready_out;
						// Trace: src/VX_mem_switch.sv:62:5
						genvar _gv_i_111;
						for (_gv_i_111 = 0; _gv_i_111 < NUM_OUTPUTS; _gv_i_111 = _gv_i_111 + 1) begin : g_rsp_data_in
							localparam i = _gv_i_111;
							// Trace: src/VX_mem_switch.sv:63:9
							assign rsp_valid_in[i] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_valid;
							// Trace: src/VX_mem_switch.sv:64:9
							assign rsp_data_in[i * 519+:519] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_data;
							// Trace: src/VX_mem_switch.sv:65:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
						end
						// Trace: src/VX_mem_switch.sv:67:5
						VX_stream_arb #(
							.NUM_INPUTS(NUM_OUTPUTS),
							.NUM_OUTPUTS(NUM_INPUTS),
							.DATAW(RSP_DATAW),
							.ARBITER(ARBITER),
							.OUT_BUF(RSP_OUT_BUF)
						) rsp_arb(
							.clk(clk),
							.reset(reset),
							.valid_in(rsp_valid_in),
							.data_in(rsp_data_in),
							.ready_in(rsp_ready_in),
							.valid_out(rsp_valid_out),
							.data_out(rsp_data_out),
							.ready_out(rsp_ready_out),
							.sel_out()
						);
						// Trace: src/VX_mem_switch.sv:84:5
						genvar _gv_i_112;
						for (_gv_i_112 = 0; _gv_i_112 < NUM_INPUTS; _gv_i_112 = _gv_i_112 + 1) begin : g_rsp_data_out
							localparam i = _gv_i_112;
							// Trace: src/VX_mem_switch.sv:85:9
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
							// Trace: src/VX_mem_switch.sv:86:9
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 519+:519];
							// Trace: src/VX_mem_switch.sv:87:9
							assign rsp_ready_out[i] = Vortex.per_cluster_mem_bus_if[i + _mbase_bus_in_if].rsp_ready;
						end
					end
					assign core_bus_nc_switch.clk = clk;
					assign core_bus_nc_switch.reset = reset;
					assign core_bus_nc_switch.bus_sel = core_req_nc_sel;
					// Trace: src/VX_cache_bypass.sv:58:5
					// expanded interface instance: core_bus_in_nc_if
					localparam _param_C0263_DATA_SIZE = WORD_SIZE;
					localparam _param_C0263_TAG_WIDTH = CORE_TAG_WIDTH;
					genvar _arr_C0263;
					for (_arr_C0263 = 0; _arr_C0263 <= 0; _arr_C0263 = _arr_C0263 + 1) begin : core_bus_in_nc_if
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_C0263_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
						localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
						localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_C0263_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:8:5
						localparam VX_gpu_pkg_UUID_WIDTH = 1;
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:12:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:20:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:24:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire [612:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire [518:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:30:5
						// Trace: src/VX_mem_bus_if.sv:38:5
					end
					// Trace: src/VX_cache_bypass.sv:62:5
					genvar _gv_i_57;
					for (_gv_i_57 = 0; _gv_i_57 < NUM_REQS; _gv_i_57 = _gv_i_57 + 1) begin : g_core_bus_nc_switch_if
						localparam i = _gv_i_57;
						// Trace: src/VX_cache_bypass.sv:63:9
						assign core_bus_in_nc_if[i].req_valid = core_bus_nc_switch_if[0 + i].req_valid;
						// Trace: src/VX_cache_bypass.sv:64:9
						assign core_bus_in_nc_if[i].req_data = core_bus_nc_switch_if[0 + i].req_data;
						// Trace: src/VX_cache_bypass.sv:65:9
						assign core_bus_nc_switch_if[0 + i].req_ready = core_bus_in_nc_if[i].req_ready;
						// Trace: src/VX_cache_bypass.sv:66:9
						assign core_bus_nc_switch_if[0 + i].rsp_valid = core_bus_in_nc_if[i].rsp_valid;
						// Trace: src/VX_cache_bypass.sv:67:9
						assign core_bus_nc_switch_if[0 + i].rsp_data = core_bus_in_nc_if[i].rsp_data;
						// Trace: src/VX_cache_bypass.sv:68:9
						assign core_bus_in_nc_if[i].rsp_ready = core_bus_nc_switch_if[0 + i].rsp_ready;
						if (CACHE_ENABLE) begin : g_cache
							// Trace: src/VX_cache_bypass.sv:70:13
							assign Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = core_bus_nc_switch_if[1 + i].req_valid;
							// Trace: src/VX_cache_bypass.sv:71:13
							assign Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = core_bus_nc_switch_if[1 + i].req_data;
							// Trace: src/VX_cache_bypass.sv:72:13
							assign core_bus_nc_switch_if[1 + i].req_ready = Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_ready;
							// Trace: src/VX_cache_bypass.sv:73:13
							assign core_bus_nc_switch_if[1 + i].rsp_valid = Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_valid;
							// Trace: src/VX_cache_bypass.sv:74:13
							assign core_bus_nc_switch_if[1 + i].rsp_data = Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_data;
							// Trace: src/VX_cache_bypass.sv:75:13
							assign Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = core_bus_nc_switch_if[1 + i].rsp_ready;
						end
						else begin : g_no_cache
							// Trace: src/VX_cache_bypass.sv:77:5
							assign Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = 0;
							// Trace: src/VX_cache_bypass.sv:78:5
							assign Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = 1'sb0;
							// Trace: src/VX_cache_bypass.sv:79:5
							assign Vortex.l3cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = 0;
						end
					end
					// Trace: src/VX_cache_bypass.sv:82:5
					// expanded interface instance: core_bus_nc_arb_if
					localparam _param_D50AC_DATA_SIZE = WORD_SIZE;
					localparam _param_D50AC_TAG_WIDTH = MEM_TAG_NC1_WIDTH;
					genvar _arr_D50AC;
					for (_arr_D50AC = 0; _arr_D50AC <= 0; _arr_D50AC = _arr_D50AC + 1) begin : core_bus_nc_arb_if
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_D50AC_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
						localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
						localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_D50AC_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:8:5
						localparam VX_gpu_pkg_UUID_WIDTH = 1;
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:12:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:20:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:24:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire [612:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire [518:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:30:5
						// Trace: src/VX_mem_bus_if.sv:38:5
					end
					// Trace: src/VX_cache_bypass.sv:86:5
					// expanded module instance: core_bus_nc_arb
					localparam _bbase_1376F_bus_in_if = 0;
					localparam _bbase_1376F_bus_out_if = 0;
					localparam _param_1376F_NUM_INPUTS = NUM_REQS;
					localparam _param_1376F_NUM_OUTPUTS = MEM_PORTS;
					localparam _param_1376F_DATA_SIZE = WORD_SIZE;
					localparam _param_1376F_TAG_WIDTH = CORE_TAG_WIDTH;
					localparam _param_1376F_TAG_SEL_IDX = TAG_SEL_IDX;
					localparam _param_1376F_ARBITER = (CACHE_ENABLE ? "P" : "R");
					localparam _param_1376F_REQ_OUT_BUF = 0;
					localparam _param_1376F_RSP_OUT_BUF = 0;
					if (1) begin : core_bus_nc_arb
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_mem_arb.sv:2:15
						localparam NUM_INPUTS = _param_1376F_NUM_INPUTS;
						// Trace: src/VX_mem_arb.sv:3:15
						localparam NUM_OUTPUTS = _param_1376F_NUM_OUTPUTS;
						// Trace: src/VX_mem_arb.sv:4:15
						localparam DATA_SIZE = _param_1376F_DATA_SIZE;
						// Trace: src/VX_mem_arb.sv:5:15
						localparam TAG_WIDTH = _param_1376F_TAG_WIDTH;
						// Trace: src/VX_mem_arb.sv:6:15
						localparam TAG_SEL_IDX = _param_1376F_TAG_SEL_IDX;
						// Trace: src/VX_mem_arb.sv:7:15
						localparam REQ_OUT_BUF = _param_1376F_REQ_OUT_BUF;
						// Trace: src/VX_mem_arb.sv:8:15
						localparam RSP_OUT_BUF = _param_1376F_RSP_OUT_BUF;
						// Trace: src/VX_mem_arb.sv:9:15
						localparam ARBITER = _param_1376F_ARBITER;
						// Trace: src/VX_mem_arb.sv:10:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_arb.sv:11:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_arb.sv:12:15
						localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
						localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
						localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
						// Trace: src/VX_mem_arb.sv:14:5
						wire clk;
						// Trace: src/VX_mem_arb.sv:15:5
						wire reset;
						// Trace: src/VX_mem_arb.sv:16:5
						localparam _mbase_bus_in_if = 0;
						// Trace: src/VX_mem_arb.sv:17:5
						localparam _mbase_bus_out_if = 0;
						// Trace: src/VX_mem_arb.sv:19:5
						localparam DATA_WIDTH = 512;
						// Trace: src/VX_mem_arb.sv:20:5
						localparam LOG_NUM_REQS = 0;
						// Trace: src/VX_mem_arb.sv:21:5
						localparam REQ_DATAW = 613;
						// Trace: src/VX_mem_arb.sv:22:5
						localparam RSP_DATAW = 519;
						// Trace: src/VX_mem_arb.sv:23:5
						localparam SEL_COUNT = NUM_OUTPUTS;
						// Trace: src/VX_mem_arb.sv:24:5
						wire [0:0] req_valid_in;
						// Trace: src/VX_mem_arb.sv:25:5
						wire [612:0] req_data_in;
						// Trace: src/VX_mem_arb.sv:26:5
						wire [0:0] req_ready_in;
						// Trace: src/VX_mem_arb.sv:27:5
						wire [0:0] req_valid_out;
						// Trace: src/VX_mem_arb.sv:28:5
						wire [612:0] req_data_out;
						// Trace: src/VX_mem_arb.sv:29:5
						wire [0:0] req_sel_out;
						// Trace: src/VX_mem_arb.sv:30:5
						wire [0:0] req_ready_out;
						// Trace: src/VX_mem_arb.sv:31:5
						genvar _gv_i_183;
						for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
							localparam i = _gv_i_183;
							// Trace: src/VX_mem_arb.sv:32:9
							assign req_valid_in[i] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_valid;
							// Trace: src/VX_mem_arb.sv:33:9
							assign req_data_in[i * 613+:613] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_data;
							// Trace: src/VX_mem_arb.sv:34:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
						end
						// Trace: src/VX_mem_arb.sv:36:5
						VX_stream_arb #(
							.NUM_INPUTS(NUM_INPUTS),
							.NUM_OUTPUTS(NUM_OUTPUTS),
							.DATAW(REQ_DATAW),
							.ARBITER(ARBITER),
							.OUT_BUF(REQ_OUT_BUF)
						) req_arb(
							.clk(clk),
							.reset(reset),
							.valid_in(req_valid_in),
							.ready_in(req_ready_in),
							.data_in(req_data_in),
							.data_out(req_data_out),
							.sel_out(req_sel_out),
							.valid_out(req_valid_out),
							.ready_out(req_ready_out)
						);
						// Trace: src/VX_mem_arb.sv:53:5
						genvar _gv_i_184;
						for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
							localparam i = _gv_i_184;
							// Trace: src/VX_mem_arb.sv:54:9
							wire [6:0] req_tag_out;
							// Trace: src/VX_mem_arb.sv:55:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
							// Trace: src/VX_mem_arb.sv:56:9
							assign {Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[612], Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[611-:26], Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[585-:512], Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[73-:64], Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[9-:3], req_tag_out} = req_data_out[i * 613+:613];
							// Trace: src/VX_mem_arb.sv:64:9
							assign req_ready_out[i] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_ready;
							if (1) begin : g_req_tag_out
								// Trace: src/VX_mem_arb.sv:76:13
								assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[6-:7] = req_tag_out;
							end
						end
						// Trace: src/VX_mem_arb.sv:79:5
						wire [0:0] rsp_valid_out;
						// Trace: src/VX_mem_arb.sv:80:5
						wire [518:0] rsp_data_out;
						// Trace: src/VX_mem_arb.sv:81:5
						wire [0:0] rsp_ready_out;
						// Trace: src/VX_mem_arb.sv:82:5
						wire [0:0] rsp_valid_in;
						// Trace: src/VX_mem_arb.sv:83:5
						wire [518:0] rsp_data_in;
						// Trace: src/VX_mem_arb.sv:84:5
						wire [0:0] rsp_ready_in;
						// Trace: src/VX_mem_arb.sv:85:5
						if (1) begin : g_rsp_arb
							genvar _gv_i_186;
							for (_gv_i_186 = 0; _gv_i_186 < NUM_OUTPUTS; _gv_i_186 = _gv_i_186 + 1) begin : g_rsp_data_in
								localparam i = _gv_i_186;
								// Trace: src/VX_mem_arb.sv:120:13
								assign rsp_valid_in[i] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_valid;
								// Trace: src/VX_mem_arb.sv:121:13
								assign rsp_data_in[i * 519+:519] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_data;
								// Trace: src/VX_mem_arb.sv:122:13
								assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
							end
							// Trace: src/VX_mem_arb.sv:124:9
							VX_stream_arb #(
								.NUM_INPUTS(NUM_OUTPUTS),
								.NUM_OUTPUTS(NUM_INPUTS),
								.DATAW(RSP_DATAW),
								.ARBITER(ARBITER),
								.OUT_BUF(RSP_OUT_BUF)
							) req_arb(
								.clk(clk),
								.reset(reset),
								.valid_in(rsp_valid_in),
								.ready_in(rsp_ready_in),
								.data_in(rsp_data_in),
								.data_out(rsp_data_out),
								.valid_out(rsp_valid_out),
								.ready_out(rsp_ready_out),
								.sel_out()
							);
						end
						// Trace: src/VX_mem_arb.sv:142:5
						genvar _gv_i_187;
						for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
							localparam i = _gv_i_187;
							// Trace: src/VX_mem_arb.sv:143:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
							// Trace: src/VX_mem_arb.sv:144:9
							assign Vortex.l3cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 519+:519];
							// Trace: src/VX_mem_arb.sv:145:9
							assign rsp_ready_out[i] = Vortex.l3cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_ready;
						end
					end
					assign core_bus_nc_arb.clk = clk;
					assign core_bus_nc_arb.reset = reset;
					// Trace: src/VX_cache_bypass.sv:101:5
					// expanded interface instance: mem_bus_out_nc_if
					localparam _param_0061C_DATA_SIZE = LINE_SIZE;
					localparam _param_0061C_TAG_WIDTH = MEM_TAG_NC2_WIDTH;
					genvar _arr_0061C;
					for (_arr_0061C = 0; _arr_0061C <= 0; _arr_0061C = _arr_0061C + 1) begin : mem_bus_out_nc_if
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_0061C_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
						localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
						localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_0061C_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:8:5
						localparam VX_gpu_pkg_UUID_WIDTH = 1;
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:12:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:20:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:24:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire [612:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire [518:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:30:5
						// Trace: src/VX_mem_bus_if.sv:38:5
					end
					// Trace: src/VX_cache_bypass.sv:105:5
					genvar _gv_i_58;
					localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
					localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
					for (_gv_i_58 = 0; _gv_i_58 < MEM_PORTS; _gv_i_58 = _gv_i_58 + 1) begin : g_mem_bus_out_nc
						localparam i = _gv_i_58;
						// Trace: src/VX_cache_bypass.sv:106:9
						wire core_req_nc_arb_rw;
						// Trace: src/VX_cache_bypass.sv:107:9
						wire [63:0] core_req_nc_arb_byteen;
						// Trace: src/VX_cache_bypass.sv:108:9
						wire [25:0] core_req_nc_arb_addr;
						// Trace: src/VX_cache_bypass.sv:109:9
						wire [2:0] core_req_nc_arb_flags;
						// Trace: src/VX_cache_bypass.sv:110:9
						wire [511:0] core_req_nc_arb_data;
						// Trace: src/VX_cache_bypass.sv:111:9
						wire [6:0] core_req_nc_arb_tag;
						// Trace: src/VX_cache_bypass.sv:112:9
						assign {core_req_nc_arb_rw, core_req_nc_arb_addr, core_req_nc_arb_data, core_req_nc_arb_byteen, core_req_nc_arb_flags, core_req_nc_arb_tag} = core_bus_nc_arb_if[i].req_data;
						// Trace: src/VX_cache_bypass.sv:120:9
						wire [25:0] core_req_nc_arb_addr_w;
						// Trace: src/VX_cache_bypass.sv:121:9
						wire [63:0] core_req_nc_arb_byteen_w;
						// Trace: src/VX_cache_bypass.sv:122:9
						wire [511:0] core_req_nc_arb_data_w;
						// Trace: src/VX_cache_bypass.sv:123:9
						wire [511:0] core_rsp_nc_arb_data_w;
						// Trace: src/VX_cache_bypass.sv:124:9
						wire [6:0] core_req_nc_arb_tag_w;
						// Trace: src/VX_cache_bypass.sv:125:9
						wire [6:0] core_rsp_nc_arb_tag_w;
						if (1) begin : g_single_word_line
							// Trace: src/VX_cache_bypass.sv:156:13
							assign core_req_nc_arb_addr_w = core_req_nc_arb_addr;
							// Trace: src/VX_cache_bypass.sv:157:13
							assign core_req_nc_arb_byteen_w = core_req_nc_arb_byteen;
							// Trace: src/VX_cache_bypass.sv:158:13
							assign core_req_nc_arb_data_w = core_req_nc_arb_data;
							// Trace: src/VX_cache_bypass.sv:159:13
							assign core_req_nc_arb_tag_w = core_req_nc_arb_tag;
							// Trace: src/VX_cache_bypass.sv:160:13
							assign core_rsp_nc_arb_data_w = mem_bus_out_nc_if[i].rsp_data[518-:512];
							// Trace: src/VX_cache_bypass.sv:161:13
							assign core_rsp_nc_arb_tag_w = sv2v_cast_7(mem_bus_out_nc_if[i].rsp_data[6-:7]);
						end
						// Trace: src/VX_cache_bypass.sv:163:9
						assign mem_bus_out_nc_if[i].req_valid = core_bus_nc_arb_if[i].req_valid;
						// Trace: src/VX_cache_bypass.sv:164:9
						assign mem_bus_out_nc_if[i].req_data = {core_req_nc_arb_rw, core_req_nc_arb_addr_w, core_req_nc_arb_data_w, core_req_nc_arb_byteen_w, core_req_nc_arb_flags, core_req_nc_arb_tag_w};
						// Trace: src/VX_cache_bypass.sv:172:9
						assign core_bus_nc_arb_if[i].req_ready = mem_bus_out_nc_if[i].req_ready;
						// Trace: src/VX_cache_bypass.sv:173:9
						assign core_bus_nc_arb_if[i].rsp_valid = mem_bus_out_nc_if[i].rsp_valid;
						// Trace: src/VX_cache_bypass.sv:174:9
						assign core_bus_nc_arb_if[i].rsp_data = {core_rsp_nc_arb_data_w, core_rsp_nc_arb_tag_w};
						// Trace: src/VX_cache_bypass.sv:178:9
						assign mem_bus_out_nc_if[i].rsp_ready = core_bus_nc_arb_if[i].rsp_ready;
					end
					// Trace: src/VX_cache_bypass.sv:180:5
					// expanded interface instance: mem_bus_out_src_if
					localparam _param_913F6_DATA_SIZE = LINE_SIZE;
					localparam _param_913F6_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
					genvar _arr_913F6;
					for (_arr_913F6 = 0; _arr_913F6 <= (((CACHE_ENABLE ? 2 : 1) * MEM_PORTS) - 1); _arr_913F6 = _arr_913F6 + 1) begin : mem_bus_out_src_if
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_913F6_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
						localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
						localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_913F6_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:8:5
						localparam VX_gpu_pkg_UUID_WIDTH = 1;
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:12:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:20:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:24:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire [(606 + (_param_913F6_TAG_WIDTH + 0)) - 1:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire [(512 + (_param_913F6_TAG_WIDTH + 0)) - 1:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:30:5
						// Trace: src/VX_mem_bus_if.sv:38:5
					end
					// Trace: src/VX_cache_bypass.sv:184:5
					genvar _gv_i_59;
					for (_gv_i_59 = 0; _gv_i_59 < MEM_PORTS; _gv_i_59 = _gv_i_59 + 1) begin : g_mem_bus_out_src
						localparam i = _gv_i_59;
						// Trace: src/VX_cache_bypass.sv:186:5
						assign mem_bus_out_src_if[0 + i].req_valid = mem_bus_out_nc_if[i].req_valid;
						// Trace: src/VX_cache_bypass.sv:187:5
						assign mem_bus_out_src_if[0 + i].req_data[539 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))] = mem_bus_out_nc_if[i].req_data[612];
						// Trace: src/VX_cache_bypass.sv:188:5
						assign mem_bus_out_src_if[0 + i].req_data[538 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))-:((602 + (_param_913F6_TAG_WIDTH + 2)) >= (579 + (_param_913F6_TAG_WIDTH + 0)) ? ((538 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))) - (512 + (_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0))))) + 1 : ((512 + (_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0)))) - (538 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)))) + 1)] = mem_bus_out_nc_if[i].req_data[611-:26];
						// Trace: src/VX_cache_bypass.sv:189:5
						assign mem_bus_out_src_if[0 + i].req_data[512 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))-:((576 + (_param_913F6_TAG_WIDTH + 2)) >= (67 + (_param_913F6_TAG_WIDTH + 0)) ? ((512 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))) - (_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0)))) + 1 : ((_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0))) - (512 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)))) + 1)] = mem_bus_out_nc_if[i].req_data[585-:512];
						// Trace: src/VX_cache_bypass.sv:190:5
						assign mem_bus_out_src_if[0 + i].req_data[_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)-:((64 + (_param_913F6_TAG_WIDTH + 2)) >= (3 + (_param_913F6_TAG_WIDTH + 0)) ? ((_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)) - (3 + (_param_913F6_TAG_WIDTH + 0))) + 1 : ((3 + (_param_913F6_TAG_WIDTH + 0)) - (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))) + 1)] = mem_bus_out_nc_if[i].req_data[73-:64];
						// Trace: src/VX_cache_bypass.sv:191:5
						assign mem_bus_out_src_if[0 + i].req_data[_param_913F6_TAG_WIDTH + 2-:((_param_913F6_TAG_WIDTH + 2) >= (_param_913F6_TAG_WIDTH + 0) ? ((_param_913F6_TAG_WIDTH + 2) - (_param_913F6_TAG_WIDTH + 0)) + 1 : ((_param_913F6_TAG_WIDTH + 0) - (_param_913F6_TAG_WIDTH + 2)) + 1)] = mem_bus_out_nc_if[i].req_data[9-:3];
						if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk1
							if (1) begin : genblk1
								if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
									// Trace: src/VX_cache_bypass.sv:195:17
									assign mem_bus_out_src_if[0 + i].req_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0] = {mem_bus_out_nc_if[i].req_data[6-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_NC2_WIDTH {1'b0}}, mem_bus_out_nc_if[i].req_data[5-:6]};
								end
								else begin : genblk1
									// Trace: src/VX_cache_bypass.sv:197:17
									assign mem_bus_out_src_if[0 + i].req_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0] = {mem_bus_out_nc_if[i].req_data[6-:1], mem_bus_out_nc_if[i].req_data[6 - (1 + (6 - (MEM_TAG_OUT_WIDTH - VX_gpu_pkg_UUID_WIDTH))):0]};
								end
							end
						end
						else begin : genblk1
							// Trace: src/VX_cache_bypass.sv:207:9
							assign mem_bus_out_src_if[0 + i].req_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0] = mem_bus_out_nc_if[i].req_data[6-:7];
						end
						// Trace: src/VX_cache_bypass.sv:209:5
						assign mem_bus_out_nc_if[i].req_ready = mem_bus_out_src_if[0 + i].req_ready;
						// Trace: src/VX_cache_bypass.sv:210:5
						assign mem_bus_out_nc_if[i].rsp_valid = mem_bus_out_src_if[0 + i].rsp_valid;
						// Trace: src/VX_cache_bypass.sv:211:5
						assign mem_bus_out_nc_if[i].rsp_data[518-:512] = mem_bus_out_src_if[0 + i].rsp_data[_param_913F6_TAG_WIDTH + 511-:((_param_913F6_TAG_WIDTH + 511) >= (_param_913F6_TAG_WIDTH + 0) ? ((_param_913F6_TAG_WIDTH + 511) - (_param_913F6_TAG_WIDTH + 0)) + 1 : ((_param_913F6_TAG_WIDTH + 0) - (_param_913F6_TAG_WIDTH + 511)) + 1)];
						if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk2
							if (1) begin : genblk1
								if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
									// Trace: src/VX_cache_bypass.sv:215:17
									assign mem_bus_out_nc_if[i].rsp_data[6-:7] = {mem_bus_out_src_if[0 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1))-:((_param_913F6_TAG_WIDTH - 1) >= (_param_913F6_TAG_WIDTH - 1) ? ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1 : ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1)], mem_bus_out_src_if[0 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 2) - (_param_913F6_TAG_WIDTH - 7))):(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 2) - (_param_913F6_TAG_WIDTH - 2)))]};
								end
								else begin : genblk1
									// Trace: src/VX_cache_bypass.sv:217:17
									assign mem_bus_out_nc_if[i].rsp_data[6-:7] = {mem_bus_out_src_if[0 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1))-:((_param_913F6_TAG_WIDTH - 1) >= (_param_913F6_TAG_WIDTH - 1) ? ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1 : ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1)], {MEM_TAG_NC2_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[0 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 2))-:_param_913F6_TAG_WIDTH - 1]};
								end
							end
						end
						else begin : genblk2
							// Trace: src/VX_cache_bypass.sv:227:9
							assign mem_bus_out_nc_if[i].rsp_data[6-:7] = mem_bus_out_src_if[0 + i].rsp_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0];
						end
						// Trace: src/VX_cache_bypass.sv:229:5
						assign mem_bus_out_src_if[0 + i].rsp_ready = mem_bus_out_nc_if[i].rsp_ready;
						if (CACHE_ENABLE) begin : g_cache
							// Trace: src/VX_cache_bypass.sv:233:5
							assign mem_bus_out_src_if[1 + i].req_valid = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_valid;
							// Trace: src/VX_cache_bypass.sv:234:5
							assign mem_bus_out_src_if[1 + i].req_data[539 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))] = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[610];
							// Trace: src/VX_cache_bypass.sv:235:5
							assign mem_bus_out_src_if[1 + i].req_data[538 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))-:((602 + (_param_913F6_TAG_WIDTH + 2)) >= (579 + (_param_913F6_TAG_WIDTH + 0)) ? ((538 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))) - (512 + (_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0))))) + 1 : ((512 + (_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0)))) - (538 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)))) + 1)] = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[609-:26];
							// Trace: src/VX_cache_bypass.sv:236:5
							assign mem_bus_out_src_if[1 + i].req_data[512 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))-:((576 + (_param_913F6_TAG_WIDTH + 2)) >= (67 + (_param_913F6_TAG_WIDTH + 0)) ? ((512 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))) - (_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0)))) + 1 : ((_param_913F6_DATA_SIZE + (3 + (_param_913F6_TAG_WIDTH + 0))) - (512 + (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)))) + 1)] = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[583-:512];
							// Trace: src/VX_cache_bypass.sv:237:5
							assign mem_bus_out_src_if[1 + i].req_data[_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)-:((64 + (_param_913F6_TAG_WIDTH + 2)) >= (3 + (_param_913F6_TAG_WIDTH + 0)) ? ((_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2)) - (3 + (_param_913F6_TAG_WIDTH + 0))) + 1 : ((3 + (_param_913F6_TAG_WIDTH + 0)) - (_param_913F6_DATA_SIZE + (_param_913F6_TAG_WIDTH + 2))) + 1)] = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[71-:64];
							// Trace: src/VX_cache_bypass.sv:238:5
							assign mem_bus_out_src_if[1 + i].req_data[_param_913F6_TAG_WIDTH + 2-:((_param_913F6_TAG_WIDTH + 2) >= (_param_913F6_TAG_WIDTH + 0) ? ((_param_913F6_TAG_WIDTH + 2) - (_param_913F6_TAG_WIDTH + 0)) + 1 : ((_param_913F6_TAG_WIDTH + 0) - (_param_913F6_TAG_WIDTH + 2)) + 1)] = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[7-:3];
							if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk1
								if (1) begin : genblk1
									if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
										// Trace: src/VX_cache_bypass.sv:242:17
										assign mem_bus_out_src_if[1 + i].req_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0] = {Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_IN_WIDTH {1'b0}}, Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[3-:4]};
									end
									else begin : genblk1
										// Trace: src/VX_cache_bypass.sv:244:17
										assign mem_bus_out_src_if[1 + i].req_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0] = {Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4 - (1 + (4 - (MEM_TAG_OUT_WIDTH - VX_gpu_pkg_UUID_WIDTH))):0]};
									end
								end
							end
							else begin : genblk1
								// Trace: src/VX_cache_bypass.sv:254:9
								assign mem_bus_out_src_if[1 + i].req_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0] = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:5];
							end
							// Trace: src/VX_cache_bypass.sv:256:5
							assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = mem_bus_out_src_if[1 + i].req_ready;
							// Trace: src/VX_cache_bypass.sv:257:5
							assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = mem_bus_out_src_if[1 + i].rsp_valid;
							// Trace: src/VX_cache_bypass.sv:258:5
							assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[516-:512] = mem_bus_out_src_if[1 + i].rsp_data[_param_913F6_TAG_WIDTH + 511-:((_param_913F6_TAG_WIDTH + 511) >= (_param_913F6_TAG_WIDTH + 0) ? ((_param_913F6_TAG_WIDTH + 511) - (_param_913F6_TAG_WIDTH + 0)) + 1 : ((_param_913F6_TAG_WIDTH + 0) - (_param_913F6_TAG_WIDTH + 511)) + 1)];
							if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk2
								if (1) begin : genblk1
									if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
										// Trace: src/VX_cache_bypass.sv:262:17
										assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1))-:((_param_913F6_TAG_WIDTH - 1) >= (_param_913F6_TAG_WIDTH - 1) ? ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1 : ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1)], mem_bus_out_src_if[1 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 2) - (_param_913F6_TAG_WIDTH - 5))):(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 2) - (_param_913F6_TAG_WIDTH - 2)))]};
									end
									else begin : genblk1
										// Trace: src/VX_cache_bypass.sv:264:17
										assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1))-:((_param_913F6_TAG_WIDTH - 1) >= (_param_913F6_TAG_WIDTH - 1) ? ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1 : ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 1)) + 1)], {MEM_TAG_IN_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[1 + i].rsp_data[(_param_913F6_TAG_WIDTH - 1) - ((_param_913F6_TAG_WIDTH - 1) - (_param_913F6_TAG_WIDTH - 2))-:_param_913F6_TAG_WIDTH - 1]};
									end
								end
							end
							else begin : genblk2
								// Trace: src/VX_cache_bypass.sv:274:9
								assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = mem_bus_out_src_if[1 + i].rsp_data[_param_913F6_TAG_WIDTH - 1-:_param_913F6_TAG_WIDTH + 0];
							end
							// Trace: src/VX_cache_bypass.sv:276:5
							assign mem_bus_out_src_if[1 + i].rsp_ready = Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_ready;
						end
						else begin : g_no_cache
							// Trace: src/VX_cache_bypass.sv:279:5
							assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = 0;
							// Trace: src/VX_cache_bypass.sv:280:5
							assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = 0;
							// Trace: src/VX_cache_bypass.sv:281:5
							assign Vortex.l3cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data = 1'sb0;
						end
					end
					// Trace: src/VX_cache_bypass.sv:284:5
					// expanded module instance: mem_bus_out_arb
					localparam _bbase_B06D0_bus_in_if = 0;
					localparam _bbase_B06D0_bus_out_if = 0;
					localparam _param_B06D0_NUM_INPUTS = (CACHE_ENABLE ? 2 : 1) * MEM_PORTS;
					localparam _param_B06D0_NUM_OUTPUTS = MEM_PORTS;
					localparam _param_B06D0_DATA_SIZE = LINE_SIZE;
					localparam _param_B06D0_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
					localparam _param_B06D0_ARBITER = "R";
					localparam _param_B06D0_REQ_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
					localparam _param_B06D0_RSP_OUT_BUF = 0;
					if (1) begin : mem_bus_out_arb
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_mem_arb.sv:2:15
						localparam NUM_INPUTS = _param_B06D0_NUM_INPUTS;
						// Trace: src/VX_mem_arb.sv:3:15
						localparam NUM_OUTPUTS = _param_B06D0_NUM_OUTPUTS;
						// Trace: src/VX_mem_arb.sv:4:15
						localparam DATA_SIZE = _param_B06D0_DATA_SIZE;
						// Trace: src/VX_mem_arb.sv:5:15
						localparam TAG_WIDTH = _param_B06D0_TAG_WIDTH;
						// Trace: src/VX_mem_arb.sv:6:15
						localparam TAG_SEL_IDX = 0;
						// Trace: src/VX_mem_arb.sv:7:15
						localparam REQ_OUT_BUF = _param_B06D0_REQ_OUT_BUF;
						// Trace: src/VX_mem_arb.sv:8:15
						localparam RSP_OUT_BUF = _param_B06D0_RSP_OUT_BUF;
						// Trace: src/VX_mem_arb.sv:9:15
						localparam ARBITER = _param_B06D0_ARBITER;
						// Trace: src/VX_mem_arb.sv:10:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_arb.sv:11:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_arb.sv:12:15
						localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
						localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
						localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
						// Trace: src/VX_mem_arb.sv:14:5
						wire clk;
						// Trace: src/VX_mem_arb.sv:15:5
						wire reset;
						// Trace: src/VX_mem_arb.sv:16:5
						localparam _mbase_bus_in_if = 0;
						// Trace: src/VX_mem_arb.sv:17:5
						localparam _mbase_bus_out_if = 0;
						// Trace: src/VX_mem_arb.sv:19:5
						localparam DATA_WIDTH = 512;
						// Trace: src/VX_mem_arb.sv:20:5
						localparam LOG_NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? $clog2((NUM_INPUTS + 0) / 1) : 0);
						// Trace: src/VX_mem_arb.sv:21:5
						localparam REQ_DATAW = 606 + TAG_WIDTH;
						// Trace: src/VX_mem_arb.sv:22:5
						localparam RSP_DATAW = DATA_WIDTH + TAG_WIDTH;
						// Trace: src/VX_mem_arb.sv:23:5
						localparam SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
						// Trace: src/VX_mem_arb.sv:24:5
						wire [NUM_INPUTS - 1:0] req_valid_in;
						// Trace: src/VX_mem_arb.sv:25:5
						wire [(NUM_INPUTS * REQ_DATAW) - 1:0] req_data_in;
						// Trace: src/VX_mem_arb.sv:26:5
						wire [NUM_INPUTS - 1:0] req_ready_in;
						// Trace: src/VX_mem_arb.sv:27:5
						wire [0:0] req_valid_out;
						// Trace: src/VX_mem_arb.sv:28:5
						wire [REQ_DATAW - 1:0] req_data_out;
						// Trace: src/VX_mem_arb.sv:29:5
						wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] req_sel_out;
						// Trace: src/VX_mem_arb.sv:30:5
						wire [0:0] req_ready_out;
						// Trace: src/VX_mem_arb.sv:31:5
						genvar _gv_i_183;
						for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
							localparam i = _gv_i_183;
							// Trace: src/VX_mem_arb.sv:32:9
							assign req_valid_in[i] = Vortex.l3cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_valid;
							// Trace: src/VX_mem_arb.sv:33:9
							assign req_data_in[i * REQ_DATAW+:REQ_DATAW] = Vortex.l3cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_data;
							// Trace: src/VX_mem_arb.sv:34:9
							assign Vortex.l3cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
						end
						// Trace: src/VX_mem_arb.sv:36:5
						VX_stream_arb #(
							.NUM_INPUTS(NUM_INPUTS),
							.NUM_OUTPUTS(NUM_OUTPUTS),
							.DATAW(REQ_DATAW),
							.ARBITER(ARBITER),
							.OUT_BUF(REQ_OUT_BUF)
						) req_arb(
							.clk(clk),
							.reset(reset),
							.valid_in(req_valid_in),
							.ready_in(req_ready_in),
							.data_in(req_data_in),
							.data_out(req_data_out),
							.sel_out(req_sel_out),
							.valid_out(req_valid_out),
							.ready_out(req_ready_out)
						);
						// Trace: src/VX_mem_arb.sv:53:5
						genvar _gv_i_184;
						for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
							localparam i = _gv_i_184;
							// Trace: src/VX_mem_arb.sv:54:9
							wire [TAG_WIDTH - 1:0] req_tag_out;
							// Trace: src/VX_mem_arb.sv:55:9
							assign Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
							// Trace: src/VX_mem_arb.sv:56:9
							assign {Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[539 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))], Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[538 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))-:((602 + (_param_4FE36_TAG_WIDTH + 2)) >= (579 + (_param_4FE36_TAG_WIDTH + 0)) ? ((538 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))) - (512 + (_param_4FE36_DATA_SIZE + (3 + (_param_4FE36_TAG_WIDTH + 0))))) + 1 : ((512 + (_param_4FE36_DATA_SIZE + (3 + (_param_4FE36_TAG_WIDTH + 0)))) - (538 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2)))) + 1)], Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[512 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))-:((576 + (_param_4FE36_TAG_WIDTH + 2)) >= (67 + (_param_4FE36_TAG_WIDTH + 0)) ? ((512 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))) - (_param_4FE36_DATA_SIZE + (3 + (_param_4FE36_TAG_WIDTH + 0)))) + 1 : ((_param_4FE36_DATA_SIZE + (3 + (_param_4FE36_TAG_WIDTH + 0))) - (512 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2)))) + 1)], Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2)-:((64 + (_param_4FE36_TAG_WIDTH + 2)) >= (3 + (_param_4FE36_TAG_WIDTH + 0)) ? ((_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2)) - (3 + (_param_4FE36_TAG_WIDTH + 0))) + 1 : ((3 + (_param_4FE36_TAG_WIDTH + 0)) - (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))) + 1)], Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[_param_4FE36_TAG_WIDTH + 2-:((_param_4FE36_TAG_WIDTH + 2) >= (_param_4FE36_TAG_WIDTH + 0) ? ((_param_4FE36_TAG_WIDTH + 2) - (_param_4FE36_TAG_WIDTH + 0)) + 1 : ((_param_4FE36_TAG_WIDTH + 0) - (_param_4FE36_TAG_WIDTH + 2)) + 1)], req_tag_out} = req_data_out[i * REQ_DATAW+:REQ_DATAW];
							// Trace: src/VX_mem_arb.sv:64:9
							assign req_ready_out[i] = Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
							if (NUM_INPUTS > NUM_OUTPUTS) begin : g_req_tag_sel_out
								// Trace: src/VX_mem_arb.sv:66:13
								VX_bits_insert #(
									.N(TAG_WIDTH),
									.S(LOG_NUM_REQS),
									.POS(TAG_SEL_IDX)
								) bits_insert(
									.data_in(req_tag_out),
									.ins_in(req_sel_out[i * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)+:(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)]),
									.data_out(Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[_param_4FE36_TAG_WIDTH - 1-:_param_4FE36_TAG_WIDTH + 0])
								);
							end
							else begin : g_req_tag_out
								// Trace: src/VX_mem_arb.sv:76:13
								assign Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[_param_4FE36_TAG_WIDTH - 1-:_param_4FE36_TAG_WIDTH + 0] = req_tag_out;
							end
						end
						// Trace: src/VX_mem_arb.sv:79:5
						wire [NUM_INPUTS - 1:0] rsp_valid_out;
						// Trace: src/VX_mem_arb.sv:80:5
						wire [(NUM_INPUTS * RSP_DATAW) - 1:0] rsp_data_out;
						// Trace: src/VX_mem_arb.sv:81:5
						wire [NUM_INPUTS - 1:0] rsp_ready_out;
						// Trace: src/VX_mem_arb.sv:82:5
						wire [0:0] rsp_valid_in;
						// Trace: src/VX_mem_arb.sv:83:5
						wire [RSP_DATAW - 1:0] rsp_data_in;
						// Trace: src/VX_mem_arb.sv:84:5
						wire [0:0] rsp_ready_in;
						// Trace: src/VX_mem_arb.sv:85:5
						if (NUM_INPUTS > NUM_OUTPUTS) begin : g_rsp_select
							// Trace: src/VX_mem_arb.sv:86:9
							wire [LOG_NUM_REQS - 1:0] rsp_sel_in;
							genvar _gv_i_185;
							for (_gv_i_185 = 0; _gv_i_185 < NUM_OUTPUTS; _gv_i_185 = _gv_i_185 + 1) begin : g_rsp_data_in
								localparam i = _gv_i_185;
								// Trace: src/VX_mem_arb.sv:88:13
								wire [TAG_WIDTH - 1:0] rsp_tag_out;
								// Trace: src/VX_mem_arb.sv:89:13
								VX_bits_remove #(
									.N(TAG_WIDTH + LOG_NUM_REQS),
									.S(LOG_NUM_REQS),
									.POS(TAG_SEL_IDX)
								) bits_remove(
									.data_in(Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[_param_4FE36_TAG_WIDTH - 1-:_param_4FE36_TAG_WIDTH + 0]),
									.sel_out(rsp_sel_in[i * LOG_NUM_REQS+:LOG_NUM_REQS]),
									.data_out(rsp_tag_out)
								);
								// Trace: src/VX_mem_arb.sv:98:13
								assign rsp_valid_in[i] = Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
								// Trace: src/VX_mem_arb.sv:99:13
								assign rsp_data_in[i * RSP_DATAW+:RSP_DATAW] = {Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[_param_4FE36_TAG_WIDTH + 511-:((_param_4FE36_TAG_WIDTH + 511) >= (_param_4FE36_TAG_WIDTH + 0) ? ((_param_4FE36_TAG_WIDTH + 511) - (_param_4FE36_TAG_WIDTH + 0)) + 1 : ((_param_4FE36_TAG_WIDTH + 0) - (_param_4FE36_TAG_WIDTH + 511)) + 1)], rsp_tag_out};
								// Trace: src/VX_mem_arb.sv:100:13
								assign Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
							end
							// Trace: src/VX_mem_arb.sv:102:9
							VX_stream_switch #(
								.NUM_INPUTS(NUM_OUTPUTS),
								.NUM_OUTPUTS(NUM_INPUTS),
								.DATAW(RSP_DATAW),
								.OUT_BUF(RSP_OUT_BUF)
							) rsp_switch(
								.clk(clk),
								.reset(reset),
								.sel_in(rsp_sel_in),
								.valid_in(rsp_valid_in),
								.ready_in(rsp_ready_in),
								.data_in(rsp_data_in),
								.data_out(rsp_data_out),
								.valid_out(rsp_valid_out),
								.ready_out(rsp_ready_out)
							);
						end
						else begin : g_rsp_arb
							genvar _gv_i_186;
							for (_gv_i_186 = 0; _gv_i_186 < NUM_OUTPUTS; _gv_i_186 = _gv_i_186 + 1) begin : g_rsp_data_in
								localparam i = _gv_i_186;
								// Trace: src/VX_mem_arb.sv:120:13
								assign rsp_valid_in[i] = Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
								// Trace: src/VX_mem_arb.sv:121:13
								assign rsp_data_in[i * RSP_DATAW+:RSP_DATAW] = Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
								// Trace: src/VX_mem_arb.sv:122:13
								assign Vortex.l3cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
							end
							// Trace: src/VX_mem_arb.sv:124:9
							VX_stream_arb #(
								.NUM_INPUTS(NUM_OUTPUTS),
								.NUM_OUTPUTS(NUM_INPUTS),
								.DATAW(RSP_DATAW),
								.ARBITER(ARBITER),
								.OUT_BUF(RSP_OUT_BUF)
							) req_arb(
								.clk(clk),
								.reset(reset),
								.valid_in(rsp_valid_in),
								.ready_in(rsp_ready_in),
								.data_in(rsp_data_in),
								.data_out(rsp_data_out),
								.valid_out(rsp_valid_out),
								.ready_out(rsp_ready_out),
								.sel_out()
							);
						end
						// Trace: src/VX_mem_arb.sv:142:5
						genvar _gv_i_187;
						for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
							localparam i = _gv_i_187;
							// Trace: src/VX_mem_arb.sv:143:9
							assign Vortex.l3cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
							// Trace: src/VX_mem_arb.sv:144:9
							assign Vortex.l3cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * RSP_DATAW+:RSP_DATAW];
							// Trace: src/VX_mem_arb.sv:145:9
							assign rsp_ready_out[i] = Vortex.l3cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_ready;
						end
					end
					assign mem_bus_out_arb.clk = clk;
					assign mem_bus_out_arb.reset = reset;
				end
				assign cache_bypass.clk = clk;
				assign cache_bypass.reset = reset;
			end
			else begin : g_no_bypass
				genvar _gv_i_38;
				for (_gv_i_38 = 0; _gv_i_38 < NUM_REQS; _gv_i_38 = _gv_i_38 + 1) begin : g_core_bus_cache_if
					localparam i = _gv_i_38;
					// Trace: src/VX_cache_wrap.sv:73:5
					assign core_bus_cache_if[i].req_valid = Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_if].req_valid;
					// Trace: src/VX_cache_wrap.sv:74:5
					assign core_bus_cache_if[i].req_data = Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_if].req_data;
					// Trace: src/VX_cache_wrap.sv:75:5
					assign Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_if].req_ready = core_bus_cache_if[i].req_ready;
					// Trace: src/VX_cache_wrap.sv:76:5
					assign Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_if].rsp_valid = core_bus_cache_if[i].rsp_valid;
					// Trace: src/VX_cache_wrap.sv:77:5
					assign Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_if].rsp_data = core_bus_cache_if[i].rsp_data;
					// Trace: src/VX_cache_wrap.sv:78:5
					assign core_bus_cache_if[i].rsp_ready = Vortex.per_cluster_mem_bus_if[i + _mbase_core_bus_if].rsp_ready;
				end
				genvar _gv_i_39;
				for (_gv_i_39 = 0; _gv_i_39 < MEM_PORTS; _gv_i_39 = _gv_i_39 + 1) begin : g_mem_bus_tmp_if
					localparam i = _gv_i_39;
					// Trace: src/VX_cache_wrap.sv:81:5
					assign mem_bus_tmp_if[i].req_valid = mem_bus_cache_if[i].req_valid;
					// Trace: src/VX_cache_wrap.sv:82:5
					assign mem_bus_tmp_if[i].req_data = mem_bus_cache_if[i].req_data;
					// Trace: src/VX_cache_wrap.sv:83:5
					assign mem_bus_cache_if[i].req_ready = mem_bus_tmp_if[i].req_ready;
					// Trace: src/VX_cache_wrap.sv:84:5
					assign mem_bus_cache_if[i].rsp_valid = mem_bus_tmp_if[i].rsp_valid;
					// Trace: src/VX_cache_wrap.sv:85:5
					assign mem_bus_cache_if[i].rsp_data = mem_bus_tmp_if[i].rsp_data;
					// Trace: src/VX_cache_wrap.sv:86:5
					assign mem_bus_tmp_if[i].rsp_ready = mem_bus_cache_if[i].rsp_ready;
				end
			end
			// Trace: src/VX_cache_wrap.sv:89:5
			genvar _gv_i_40;
			for (_gv_i_40 = 0; _gv_i_40 < MEM_PORTS; _gv_i_40 = _gv_i_40 + 1) begin : g_mem_bus_if
				localparam i = _gv_i_40;
				if (WRITE_ENABLE) begin : g_we
					// Trace: src/VX_cache_wrap.sv:91:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
					// Trace: src/VX_cache_wrap.sv:92:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[i].req_data;
					// Trace: src/VX_cache_wrap.sv:93:5
					assign mem_bus_tmp_if[i].req_ready = Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_ready;
					// Trace: src/VX_cache_wrap.sv:94:5
					assign mem_bus_tmp_if[i].rsp_valid = Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
					// Trace: src/VX_cache_wrap.sv:95:5
					assign mem_bus_tmp_if[i].rsp_data = Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
					// Trace: src/VX_cache_wrap.sv:96:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
				end
				else begin : g_ro
					// Trace: src/VX_cache_wrap.sv:98:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
					// Trace: src/VX_cache_wrap.sv:99:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data[612] = 0;
					// Trace: src/VX_cache_wrap.sv:100:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data[611-:26] = mem_bus_tmp_if[i].req_data[538 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))-:((602 + (_param_4FE36_TAG_WIDTH + 2)) >= (579 + (_param_4FE36_TAG_WIDTH + 0)) ? ((538 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2))) - (512 + (_param_4FE36_DATA_SIZE + (3 + (_param_4FE36_TAG_WIDTH + 0))))) + 1 : ((512 + (_param_4FE36_DATA_SIZE + (3 + (_param_4FE36_TAG_WIDTH + 0)))) - (538 + (_param_4FE36_DATA_SIZE + (_param_4FE36_TAG_WIDTH + 2)))) + 1)];
					// Trace: src/VX_cache_wrap.sv:101:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data[585-:512] = 1'sb0;
					// Trace: src/VX_cache_wrap.sv:102:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data[73-:64] = 1'sb1;
					// Trace: src/VX_cache_wrap.sv:103:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data[9-:3] = mem_bus_tmp_if[i].req_data[_param_4FE36_TAG_WIDTH + 2-:((_param_4FE36_TAG_WIDTH + 2) >= (_param_4FE36_TAG_WIDTH + 0) ? ((_param_4FE36_TAG_WIDTH + 2) - (_param_4FE36_TAG_WIDTH + 0)) + 1 : ((_param_4FE36_TAG_WIDTH + 0) - (_param_4FE36_TAG_WIDTH + 2)) + 1)];
					// Trace: src/VX_cache_wrap.sv:104:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_data[6-:7] = mem_bus_tmp_if[i].req_data[_param_4FE36_TAG_WIDTH - 1-:_param_4FE36_TAG_WIDTH + 0];
					// Trace: src/VX_cache_wrap.sv:105:5
					assign mem_bus_tmp_if[i].req_ready = Vortex.mem_bus_if[i + _mbase_mem_bus_if].req_ready;
					// Trace: src/VX_cache_wrap.sv:106:5
					assign mem_bus_tmp_if[i].rsp_valid = Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
					// Trace: src/VX_cache_wrap.sv:107:5
					assign mem_bus_tmp_if[i].rsp_data[_param_4FE36_TAG_WIDTH + 511-:((_param_4FE36_TAG_WIDTH + 511) >= (_param_4FE36_TAG_WIDTH + 0) ? ((_param_4FE36_TAG_WIDTH + 511) - (_param_4FE36_TAG_WIDTH + 0)) + 1 : ((_param_4FE36_TAG_WIDTH + 0) - (_param_4FE36_TAG_WIDTH + 511)) + 1)] = Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_data[518-:512];
					// Trace: src/VX_cache_wrap.sv:108:5
					assign mem_bus_tmp_if[i].rsp_data[_param_4FE36_TAG_WIDTH - 1-:_param_4FE36_TAG_WIDTH + 0] = Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_data[6-:7];
					// Trace: src/VX_cache_wrap.sv:109:5
					assign Vortex.mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
				end
			end
			// Trace: src/VX_cache_wrap.sv:112:5
			if (1) begin : g_passthru
				genvar _gv_i_41;
				for (_gv_i_41 = 0; _gv_i_41 < NUM_REQS; _gv_i_41 = _gv_i_41 + 1) begin : g_core_bus_cache_if
					localparam i = _gv_i_41;
					// Trace: src/VX_cache_wrap.sv:141:5
					assign core_bus_cache_if[i].req_ready = 0;
					// Trace: src/VX_cache_wrap.sv:142:5
					assign core_bus_cache_if[i].rsp_valid = 0;
					// Trace: src/VX_cache_wrap.sv:143:5
					assign core_bus_cache_if[i].rsp_data = 1'sb0;
				end
				genvar _gv_i_42;
				for (_gv_i_42 = 0; _gv_i_42 < MEM_PORTS; _gv_i_42 = _gv_i_42 + 1) begin : g_mem_bus_cache_if
					localparam i = _gv_i_42;
					// Trace: src/VX_cache_wrap.sv:146:5
					assign mem_bus_cache_if[i].req_valid = 0;
					// Trace: src/VX_cache_wrap.sv:147:5
					assign mem_bus_cache_if[i].req_data = 1'sb0;
					// Trace: src/VX_cache_wrap.sv:148:5
					assign mem_bus_cache_if[i].rsp_ready = 0;
				end
			end
		end
	endgenerate
	assign l3cache.clk = clk;
	assign l3cache.reset = l3_reset;
	// Trace: src/Vortex.sv:62:5
	genvar _gv_i_95;
	generate
		for (_gv_i_95 = 0; _gv_i_95 < VX_gpu_pkg_L3_NUM_REQS; _gv_i_95 = _gv_i_95 + 1) begin : g_mem_bus_if
			localparam i = _gv_i_95;
			// Trace: src/Vortex.sv:63:9
			assign mem_req_valid[i] = mem_bus_if[i].req_valid;
			// Trace: src/Vortex.sv:64:9
			assign mem_req_rw[i] = mem_bus_if[i].req_data[612];
			// Trace: src/Vortex.sv:65:9
			assign mem_req_byteen[i * 64+:64] = mem_bus_if[i].req_data[73-:64];
			// Trace: src/Vortex.sv:66:9
			assign mem_req_addr[i * 26+:26] = mem_bus_if[i].req_data[611-:26];
			// Trace: src/Vortex.sv:67:9
			assign mem_req_data[i * 512+:512] = mem_bus_if[i].req_data[585-:512];
			// Trace: src/Vortex.sv:68:9
			assign mem_req_tag[i * 7+:7] = mem_bus_if[i].req_data[6-:7];
			// Trace: src/Vortex.sv:69:9
			assign mem_bus_if[i].req_ready = mem_req_ready[i];
			// Trace: src/Vortex.sv:70:9
			assign mem_bus_if[i].rsp_valid = mem_rsp_valid[i];
			// Trace: src/Vortex.sv:71:9
			assign mem_bus_if[i].rsp_data[518-:512] = mem_rsp_data[i * 512+:512];
			// Trace: src/Vortex.sv:72:9
			assign mem_bus_if[i].rsp_data[6-:7] = mem_rsp_tag[i * 7+:7];
			// Trace: src/Vortex.sv:73:9
			assign mem_rsp_ready[i] = mem_bus_if[i].rsp_ready;
		end
	endgenerate
	// Trace: src/Vortex.sv:75:5
	// expanded interface instance: dcr_bus_if
	generate
		if (1) begin : dcr_bus_if
			// removed import VX_gpu_pkg::*;
			// Trace: src/VX_dcr_bus_if.sv:2:5
			wire write_valid;
			// Trace: src/VX_dcr_bus_if.sv:3:5
			localparam VX_gpu_pkg_VX_DCR_ADDR_WIDTH = 12;
			wire [11:0] write_addr;
			// Trace: src/VX_dcr_bus_if.sv:4:5
			localparam VX_gpu_pkg_VX_DCR_DATA_WIDTH = 32;
			wire [31:0] write_data;
			// Trace: src/VX_dcr_bus_if.sv:5:5
			// Trace: src/VX_dcr_bus_if.sv:10:5
		end
	endgenerate
	// Trace: src/Vortex.sv:76:5
	assign dcr_bus_if.write_valid = dcr_wr_valid;
	// Trace: src/Vortex.sv:77:5
	assign dcr_bus_if.write_addr = dcr_wr_addr;
	// Trace: src/Vortex.sv:78:5
	assign dcr_bus_if.write_data = dcr_wr_data;
	// Trace: src/Vortex.sv:79:5
	wire [0:0] per_cluster_busy;
	// Trace: src/Vortex.sv:80:5
	genvar _gv_cluster_id_1;
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	function automatic [29:0] sv2v_cast_30;
		input reg [29:0] inp;
		sv2v_cast_30 = inp;
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	function automatic signed [2:0] sv2v_cast_22555_signed;
		input reg signed [2:0] inp;
		sv2v_cast_22555_signed = inp;
	endfunction
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	function automatic signed [1:0] sv2v_cast_2_signed;
		input reg signed [1:0] inp;
		sv2v_cast_2_signed = inp;
	endfunction
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	function automatic signed [0:0] sv2v_cast_1_signed;
		input reg signed [0:0] inp;
		sv2v_cast_1_signed = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	function automatic [25:0] sv2v_cast_26;
		input reg [25:0] inp;
		sv2v_cast_26 = inp;
	endfunction
	function automatic [43:0] sv2v_cast_44;
		input reg [43:0] inp;
		sv2v_cast_44 = inp;
	endfunction
	generate
		for (_gv_cluster_id_1 = 0; _gv_cluster_id_1 < 1; _gv_cluster_id_1 = _gv_cluster_id_1 + 1) begin : g_clusters
			localparam cluster_id = _gv_cluster_id_1;
			// Trace: src/Vortex.sv:81:5
			wire [0:0] cluster_reset;
			// Trace: src/Vortex.sv:82:5
			VX_reset_relay #(
				.N(1),
				.MAX_FANOUT(0)
			) __cluster_reset(
				.clk(clk),
				.reset(reset),
				.reset_o(cluster_reset)
			);
			// Trace: src/Vortex.sv:87:9
			// expanded interface instance: cluster_dcr_bus_if
			if (1) begin : cluster_dcr_bus_if
				// removed import VX_gpu_pkg::*;
				// Trace: src/VX_dcr_bus_if.sv:2:5
				wire write_valid;
				// Trace: src/VX_dcr_bus_if.sv:3:5
				localparam VX_gpu_pkg_VX_DCR_ADDR_WIDTH = 12;
				wire [11:0] write_addr;
				// Trace: src/VX_dcr_bus_if.sv:4:5
				localparam VX_gpu_pkg_VX_DCR_DATA_WIDTH = 32;
				wire [31:0] write_data;
				// Trace: src/VX_dcr_bus_if.sv:5:5
				// Trace: src/VX_dcr_bus_if.sv:10:5
			end
			if (1) begin : genblk1
				// Trace: src/Vortex.sv:101:9
				assign {cluster_dcr_bus_if.write_valid, cluster_dcr_bus_if.write_addr, cluster_dcr_bus_if.write_data} = {dcr_bus_if.write_valid && 1'b1, dcr_bus_if.write_addr, dcr_bus_if.write_data};
			end
			// Trace: src/Vortex.sv:104:9
			// expanded module instance: cluster
			localparam _bbase_5867A_mem_bus_if = cluster_id * VX_gpu_pkg_L2_NUM_REQS;
			localparam _param_5867A_CLUSTER_ID = cluster_id;
			localparam _param_5867A_INSTANCE_ID = "";
			if (1) begin : cluster
				// removed import VX_gpu_pkg::*;
				// Trace: src/VX_cluster.sv:2:15
				localparam CLUSTER_ID = _param_5867A_CLUSTER_ID;
				// Trace: src/VX_cluster.sv:3:15
				localparam INSTANCE_ID = _param_5867A_INSTANCE_ID;
				// Trace: src/VX_cluster.sv:5:5
				wire clk;
				// Trace: src/VX_cluster.sv:6:5
				wire reset;
				// Trace: src/VX_cluster.sv:7:5
				// removed modport instance dcr_bus_if
				// Trace: src/VX_cluster.sv:8:5
				localparam VX_gpu_pkg_DCACHE_WORD_SIZE = 16;
				localparam VX_gpu_pkg_XLENB = 4;
				localparam VX_gpu_pkg_LSU_WORD_SIZE = VX_gpu_pkg_XLENB;
				localparam VX_gpu_pkg_DCACHE_CHANNELS = 1;
				localparam VX_gpu_pkg_DCACHE_NUM_REQS = 1;
				localparam VX_gpu_pkg_NUM_SOCKETS = 1;
				localparam VX_gpu_pkg_L2_NUM_REQS = 1;
				localparam _mbase_mem_bus_if = _bbase_5867A_mem_bus_if;
				// Trace: src/VX_cluster.sv:9:5
				wire busy;
				// Trace: src/VX_cluster.sv:11:5
				localparam VX_gpu_pkg_DCACHE_LINE_SIZE = 64;
				localparam VX_gpu_pkg_DCACHE_MERGED_REQS = 1;
				localparam VX_gpu_pkg_DCACHE_MEM_BATCHES = 1;
				localparam VX_gpu_pkg_DCACHE_TAG_ID_BITS = 2;
				localparam VX_gpu_pkg_UUID_WIDTH = 1;
				localparam VX_gpu_pkg_DCACHE_TAG_WIDTH = 3;
				localparam VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH = 6;
				localparam VX_gpu_pkg_ICACHE_MEM_TAG_WIDTH = 5;
				localparam VX_gpu_pkg_L1_MEM_TAG_WIDTH = VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH;
				localparam VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH = 7;
				// expanded interface instance: per_socket_mem_bus_if
				localparam _param_1BD2B_DATA_SIZE = 64;
				localparam _param_1BD2B_TAG_WIDTH = VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH;
				genvar _arr_1BD2B;
				for (_arr_1BD2B = 0; _arr_1BD2B <= 0; _arr_1BD2B = _arr_1BD2B + 1) begin : per_socket_mem_bus_if
					// removed import VX_gpu_pkg::*;
					// Trace: src/VX_mem_bus_if.sv:2:15
					localparam DATA_SIZE = _param_1BD2B_DATA_SIZE;
					// Trace: src/VX_mem_bus_if.sv:3:15
					localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
					localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
					localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
					// Trace: src/VX_mem_bus_if.sv:4:15
					localparam TAG_WIDTH = _param_1BD2B_TAG_WIDTH;
					// Trace: src/VX_mem_bus_if.sv:5:15
					localparam MEM_ADDR_WIDTH = 32;
					// Trace: src/VX_mem_bus_if.sv:6:15
					localparam ADDR_WIDTH = 26;
					// Trace: src/VX_mem_bus_if.sv:8:5
					localparam VX_gpu_pkg_UUID_WIDTH = 1;
					// removed localparam type tag_t
					// Trace: src/VX_mem_bus_if.sv:12:5
					// removed localparam type req_data_t
					// Trace: src/VX_mem_bus_if.sv:20:5
					// removed localparam type rsp_data_t
					// Trace: src/VX_mem_bus_if.sv:24:5
					wire req_valid;
					// Trace: src/VX_mem_bus_if.sv:25:5
					wire [612:0] req_data;
					// Trace: src/VX_mem_bus_if.sv:26:5
					wire req_ready;
					// Trace: src/VX_mem_bus_if.sv:27:5
					wire rsp_valid;
					// Trace: src/VX_mem_bus_if.sv:28:5
					wire [518:0] rsp_data;
					// Trace: src/VX_mem_bus_if.sv:29:5
					wire rsp_ready;
					// Trace: src/VX_mem_bus_if.sv:30:5
					// Trace: src/VX_mem_bus_if.sv:38:5
				end
				// Trace: src/VX_cluster.sv:15:5
				wire [0:0] l2_reset;
				// Trace: src/VX_cluster.sv:16:5
				VX_reset_relay #(
					.N(1),
					.MAX_FANOUT(0)
				) __l2_reset(
					.clk(clk),
					.reset(reset),
					.reset_o(l2_reset)
				);
				// Trace: src/VX_cluster.sv:21:5
				localparam VX_gpu_pkg_L2_TAG_WIDTH = VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH;
				localparam VX_gpu_pkg_L2_WORD_SIZE = 64;
				// expanded module instance: l2cache
				localparam _bbase_56EB4_core_bus_if = 0;
				localparam _bbase_56EB4_mem_bus_if = cluster_id * VX_gpu_pkg_L2_NUM_REQS;
				localparam _param_56EB4_INSTANCE_ID = "";
				localparam _param_56EB4_CACHE_SIZE = 1048576;
				localparam _param_56EB4_LINE_SIZE = 64;
				localparam _param_56EB4_NUM_BANKS = VX_gpu_pkg_L2_NUM_REQS;
				localparam _param_56EB4_NUM_WAYS = 8;
				localparam _param_56EB4_WORD_SIZE = VX_gpu_pkg_L2_WORD_SIZE;
				localparam _param_56EB4_NUM_REQS = VX_gpu_pkg_L2_NUM_REQS;
				localparam _param_56EB4_MEM_PORTS = VX_gpu_pkg_L2_NUM_REQS;
				localparam _param_56EB4_CRSQ_SIZE = 2;
				localparam _param_56EB4_MSHR_SIZE = 16;
				localparam _param_56EB4_MRSQ_SIZE = 4;
				localparam _param_56EB4_MREQ_SIZE = 4;
				localparam _param_56EB4_TAG_WIDTH = VX_gpu_pkg_L2_TAG_WIDTH;
				localparam _param_56EB4_WRITE_ENABLE = 1;
				localparam _param_56EB4_WRITEBACK = 0;
				localparam _param_56EB4_DIRTY_BYTES = 0;
				localparam _param_56EB4_REPL_POLICY = 1;
				localparam _param_56EB4_CORE_OUT_BUF = 3;
				localparam _param_56EB4_MEM_OUT_BUF = 3;
				localparam _param_56EB4_NC_ENABLE = 1;
				localparam _param_56EB4_PASSTHRU = 1'd1;
				if (1) begin : l2cache
					// removed import VX_gpu_pkg::*;
					// Trace: src/VX_cache_wrap.sv:2:15
					localparam INSTANCE_ID = _param_56EB4_INSTANCE_ID;
					// Trace: src/VX_cache_wrap.sv:3:15
					localparam TAG_SEL_IDX = 0;
					// Trace: src/VX_cache_wrap.sv:4:15
					localparam NUM_REQS = _param_56EB4_NUM_REQS;
					// Trace: src/VX_cache_wrap.sv:5:15
					localparam MEM_PORTS = _param_56EB4_MEM_PORTS;
					// Trace: src/VX_cache_wrap.sv:6:15
					localparam CACHE_SIZE = _param_56EB4_CACHE_SIZE;
					// Trace: src/VX_cache_wrap.sv:7:15
					localparam LINE_SIZE = _param_56EB4_LINE_SIZE;
					// Trace: src/VX_cache_wrap.sv:8:15
					localparam NUM_BANKS = _param_56EB4_NUM_BANKS;
					// Trace: src/VX_cache_wrap.sv:9:15
					localparam NUM_WAYS = _param_56EB4_NUM_WAYS;
					// Trace: src/VX_cache_wrap.sv:10:15
					localparam WORD_SIZE = _param_56EB4_WORD_SIZE;
					// Trace: src/VX_cache_wrap.sv:11:15
					localparam CRSQ_SIZE = _param_56EB4_CRSQ_SIZE;
					// Trace: src/VX_cache_wrap.sv:12:15
					localparam MSHR_SIZE = _param_56EB4_MSHR_SIZE;
					// Trace: src/VX_cache_wrap.sv:13:15
					localparam MRSQ_SIZE = _param_56EB4_MRSQ_SIZE;
					// Trace: src/VX_cache_wrap.sv:14:15
					localparam MREQ_SIZE = _param_56EB4_MREQ_SIZE;
					// Trace: src/VX_cache_wrap.sv:15:15
					localparam WRITE_ENABLE = _param_56EB4_WRITE_ENABLE;
					// Trace: src/VX_cache_wrap.sv:16:15
					localparam WRITEBACK = _param_56EB4_WRITEBACK;
					// Trace: src/VX_cache_wrap.sv:17:15
					localparam DIRTY_BYTES = _param_56EB4_DIRTY_BYTES;
					// Trace: src/VX_cache_wrap.sv:18:15
					localparam REPL_POLICY = _param_56EB4_REPL_POLICY;
					// Trace: src/VX_cache_wrap.sv:19:15
					localparam VX_gpu_pkg_UUID_WIDTH = 1;
					localparam TAG_WIDTH = _param_56EB4_TAG_WIDTH;
					// Trace: src/VX_cache_wrap.sv:20:15
					localparam NC_ENABLE = _param_56EB4_NC_ENABLE;
					// Trace: src/VX_cache_wrap.sv:21:15
					localparam PASSTHRU = _param_56EB4_PASSTHRU;
					// Trace: src/VX_cache_wrap.sv:22:15
					localparam CORE_OUT_BUF = _param_56EB4_CORE_OUT_BUF;
					// Trace: src/VX_cache_wrap.sv:23:15
					localparam MEM_OUT_BUF = _param_56EB4_MEM_OUT_BUF;
					// Trace: src/VX_cache_wrap.sv:25:5
					wire clk;
					// Trace: src/VX_cache_wrap.sv:26:5
					wire reset;
					// Trace: src/VX_cache_wrap.sv:27:5
					localparam _mbase_core_bus_if = 0;
					// Trace: src/VX_cache_wrap.sv:28:5
					localparam _mbase_mem_bus_if = _bbase_56EB4_mem_bus_if;
					// Trace: src/VX_cache_wrap.sv:30:5
					localparam CACHE_MEM_TAG_WIDTH = 5;
					// Trace: src/VX_cache_wrap.sv:32:5
					localparam BYPASS_TAG_WIDTH = 7;
					// Trace: src/VX_cache_wrap.sv:34:5
					localparam NC_TAG_WIDTH = 8;
					// Trace: src/VX_cache_wrap.sv:35:5
					localparam MEM_TAG_WIDTH = (PASSTHRU ? BYPASS_TAG_WIDTH : (NC_ENABLE ? NC_TAG_WIDTH : CACHE_MEM_TAG_WIDTH));
					// Trace: src/VX_cache_wrap.sv:36:5
					localparam BYPASS_ENABLE = 1'd1;
					// Trace: src/VX_cache_wrap.sv:37:5
					// expanded interface instance: core_bus_cache_if
					localparam _param_24C1C_DATA_SIZE = WORD_SIZE;
					localparam _param_24C1C_TAG_WIDTH = TAG_WIDTH;
					genvar _arr_24C1C;
					for (_arr_24C1C = 0; _arr_24C1C <= 0; _arr_24C1C = _arr_24C1C + 1) begin : core_bus_cache_if
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_24C1C_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
						localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
						localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_24C1C_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:8:5
						localparam VX_gpu_pkg_UUID_WIDTH = 1;
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:12:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:20:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:24:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire [612:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire [518:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:30:5
						// Trace: src/VX_mem_bus_if.sv:38:5
					end
					// Trace: src/VX_cache_wrap.sv:41:5
					// expanded interface instance: mem_bus_cache_if
					localparam _param_D895D_DATA_SIZE = LINE_SIZE;
					localparam _param_D895D_TAG_WIDTH = CACHE_MEM_TAG_WIDTH;
					genvar _arr_D895D;
					for (_arr_D895D = 0; _arr_D895D <= 0; _arr_D895D = _arr_D895D + 1) begin : mem_bus_cache_if
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_D895D_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
						localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
						localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_D895D_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:8:5
						localparam VX_gpu_pkg_UUID_WIDTH = 1;
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:12:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:20:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:24:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire [610:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire [516:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:30:5
						// Trace: src/VX_mem_bus_if.sv:38:5
					end
					// Trace: src/VX_cache_wrap.sv:45:5
					// expanded interface instance: mem_bus_tmp_if
					localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
					localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH;
					genvar _arr_4FE36;
					for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_mem_bus_if.sv:2:15
						localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
						// Trace: src/VX_mem_bus_if.sv:3:15
						localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
						localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
						localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:4:15
						localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
						// Trace: src/VX_mem_bus_if.sv:5:15
						localparam MEM_ADDR_WIDTH = 32;
						// Trace: src/VX_mem_bus_if.sv:6:15
						localparam ADDR_WIDTH = 26;
						// Trace: src/VX_mem_bus_if.sv:8:5
						localparam VX_gpu_pkg_UUID_WIDTH = 1;
						// removed localparam type tag_t
						// Trace: src/VX_mem_bus_if.sv:12:5
						// removed localparam type req_data_t
						// Trace: src/VX_mem_bus_if.sv:20:5
						// removed localparam type rsp_data_t
						// Trace: src/VX_mem_bus_if.sv:24:5
						wire req_valid;
						// Trace: src/VX_mem_bus_if.sv:25:5
						wire [612:0] req_data;
						// Trace: src/VX_mem_bus_if.sv:26:5
						wire req_ready;
						// Trace: src/VX_mem_bus_if.sv:27:5
						wire rsp_valid;
						// Trace: src/VX_mem_bus_if.sv:28:5
						wire [518:0] rsp_data;
						// Trace: src/VX_mem_bus_if.sv:29:5
						wire rsp_ready;
						// Trace: src/VX_mem_bus_if.sv:30:5
						// Trace: src/VX_mem_bus_if.sv:38:5
					end
					// Trace: src/VX_cache_wrap.sv:49:5
					if (BYPASS_ENABLE) begin : g_bypass
						// Trace: src/VX_cache_wrap.sv:50:9
						// expanded module instance: cache_bypass
						localparam _bbase_714AA_core_bus_in_if = 0;
						localparam _bbase_714AA_core_bus_out_if = 0;
						localparam _bbase_714AA_mem_bus_in_if = 0;
						localparam _bbase_714AA_mem_bus_out_if = 0;
						localparam _param_714AA_NUM_REQS = NUM_REQS;
						localparam _param_714AA_MEM_PORTS = MEM_PORTS;
						localparam _param_714AA_TAG_SEL_IDX = TAG_SEL_IDX;
						localparam _param_714AA_CACHE_ENABLE = !PASSTHRU;
						localparam _param_714AA_WORD_SIZE = WORD_SIZE;
						localparam _param_714AA_LINE_SIZE = LINE_SIZE;
						localparam _param_714AA_CORE_ADDR_WIDTH = 26;
						localparam _param_714AA_CORE_TAG_WIDTH = TAG_WIDTH;
						localparam _param_714AA_MEM_ADDR_WIDTH = 26;
						localparam _param_714AA_MEM_TAG_IN_WIDTH = CACHE_MEM_TAG_WIDTH;
						localparam _param_714AA_CORE_OUT_BUF = CORE_OUT_BUF;
						localparam _param_714AA_MEM_OUT_BUF = MEM_OUT_BUF;
						if (1) begin : cache_bypass
							// removed import VX_gpu_pkg::*;
							// Trace: src/VX_cache_bypass.sv:2:15
							localparam NUM_REQS = _param_714AA_NUM_REQS;
							// Trace: src/VX_cache_bypass.sv:3:15
							localparam MEM_PORTS = _param_714AA_MEM_PORTS;
							// Trace: src/VX_cache_bypass.sv:4:15
							localparam TAG_SEL_IDX = _param_714AA_TAG_SEL_IDX;
							// Trace: src/VX_cache_bypass.sv:5:15
							localparam CACHE_ENABLE = _param_714AA_CACHE_ENABLE;
							// Trace: src/VX_cache_bypass.sv:6:15
							localparam WORD_SIZE = _param_714AA_WORD_SIZE;
							// Trace: src/VX_cache_bypass.sv:7:15
							localparam LINE_SIZE = _param_714AA_LINE_SIZE;
							// Trace: src/VX_cache_bypass.sv:8:15
							localparam CORE_ADDR_WIDTH = _param_714AA_CORE_ADDR_WIDTH;
							// Trace: src/VX_cache_bypass.sv:9:15
							localparam CORE_TAG_WIDTH = _param_714AA_CORE_TAG_WIDTH;
							// Trace: src/VX_cache_bypass.sv:10:15
							localparam MEM_ADDR_WIDTH = _param_714AA_MEM_ADDR_WIDTH;
							// Trace: src/VX_cache_bypass.sv:11:15
							localparam MEM_TAG_IN_WIDTH = _param_714AA_MEM_TAG_IN_WIDTH;
							// Trace: src/VX_cache_bypass.sv:12:15
							localparam CORE_OUT_BUF = _param_714AA_CORE_OUT_BUF;
							// Trace: src/VX_cache_bypass.sv:13:15
							localparam MEM_OUT_BUF = _param_714AA_MEM_OUT_BUF;
							// Trace: src/VX_cache_bypass.sv:15:5
							wire clk;
							// Trace: src/VX_cache_bypass.sv:16:5
							wire reset;
							// Trace: src/VX_cache_bypass.sv:17:5
							localparam _mbase_core_bus_in_if = 0;
							// Trace: src/VX_cache_bypass.sv:18:5
							localparam _mbase_core_bus_out_if = 0;
							// Trace: src/VX_cache_bypass.sv:19:5
							localparam _mbase_mem_bus_in_if = 0;
							// Trace: src/VX_cache_bypass.sv:20:5
							localparam _mbase_mem_bus_out_if = 0;
							// Trace: src/VX_cache_bypass.sv:22:5
							localparam DIRECT_PASSTHRU = (!CACHE_ENABLE && 1'd1) && 1'd1;
							// Trace: src/VX_cache_bypass.sv:23:5
							localparam CORE_DATA_WIDTH = 512;
							// Trace: src/VX_cache_bypass.sv:24:5
							localparam WORDS_PER_LINE = 1;
							// Trace: src/VX_cache_bypass.sv:25:5
							localparam WSEL_BITS = 0;
							// Trace: src/VX_cache_bypass.sv:26:5
							localparam VX_gpu_pkg_UUID_WIDTH = 1;
							localparam CORE_TAG_ID_WIDTH = 6;
							// Trace: src/VX_cache_bypass.sv:27:5
							localparam MEM_TAG_ID_WIDTH = 6;
							// Trace: src/VX_cache_bypass.sv:28:5
							localparam MEM_TAG_NC1_WIDTH = 7;
							// Trace: src/VX_cache_bypass.sv:29:5
							localparam MEM_TAG_NC2_WIDTH = 7;
							// Trace: src/VX_cache_bypass.sv:30:5
							localparam MEM_TAG_OUT_WIDTH = (CACHE_ENABLE ? MEM_TAG_NC2_WIDTH : MEM_TAG_NC2_WIDTH);
							// Trace: src/VX_cache_bypass.sv:31:5
							// expanded interface instance: core_bus_nc_switch_if
							localparam _param_95306_DATA_SIZE = WORD_SIZE;
							localparam _param_95306_TAG_WIDTH = CORE_TAG_WIDTH;
							genvar _arr_95306;
							for (_arr_95306 = 0; _arr_95306 <= (((CACHE_ENABLE ? 2 : 1) * NUM_REQS) - 1); _arr_95306 = _arr_95306 + 1) begin : core_bus_nc_switch_if
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_95306_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
								localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
								localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_95306_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:8:5
								localparam VX_gpu_pkg_UUID_WIDTH = 1;
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:12:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:20:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:24:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire [612:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire [518:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:30:5
								// Trace: src/VX_mem_bus_if.sv:38:5
							end
							// Trace: src/VX_cache_bypass.sv:35:5
							wire [0:0] core_req_nc_sel;
							// Trace: src/VX_cache_bypass.sv:36:5
							genvar _gv_i_56;
							localparam VX_gpu_pkg_MEM_REQ_FLAG_IO = 1;
							for (_gv_i_56 = 0; _gv_i_56 < NUM_REQS; _gv_i_56 = _gv_i_56 + 1) begin : g_core_req_is_nc
								localparam i = _gv_i_56;
								if (CACHE_ENABLE) begin : g_cache
									// Trace: src/VX_cache_bypass.sv:38:13
									assign core_req_nc_sel[i] = ~Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_in_if].req_data[8];
								end
								else begin : g_no_cache
									// Trace: src/VX_cache_bypass.sv:40:13
									assign core_req_nc_sel[i] = 1'b0;
								end
							end
							// Trace: src/VX_cache_bypass.sv:43:5
							// expanded module instance: core_bus_nc_switch
							localparam _bbase_69FDB_bus_in_if = 0;
							localparam _bbase_69FDB_bus_out_if = 0;
							localparam _param_69FDB_NUM_INPUTS = NUM_REQS;
							localparam _param_69FDB_NUM_OUTPUTS = (CACHE_ENABLE ? 2 : 1) * NUM_REQS;
							localparam _param_69FDB_DATA_SIZE = WORD_SIZE;
							localparam _param_69FDB_TAG_WIDTH = CORE_TAG_WIDTH;
							localparam _param_69FDB_ARBITER = "R";
							localparam _param_69FDB_REQ_OUT_BUF = 0;
							localparam _param_69FDB_RSP_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
							if (1) begin : core_bus_nc_switch
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_switch.sv:2:15
								localparam NUM_INPUTS = _param_69FDB_NUM_INPUTS;
								// Trace: src/VX_mem_switch.sv:3:15
								localparam NUM_OUTPUTS = _param_69FDB_NUM_OUTPUTS;
								// Trace: src/VX_mem_switch.sv:4:15
								localparam DATA_SIZE = _param_69FDB_DATA_SIZE;
								// Trace: src/VX_mem_switch.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_switch.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_switch.sv:7:15
								localparam TAG_WIDTH = _param_69FDB_TAG_WIDTH;
								// Trace: src/VX_mem_switch.sv:8:15
								localparam REQ_OUT_BUF = _param_69FDB_REQ_OUT_BUF;
								// Trace: src/VX_mem_switch.sv:9:15
								localparam RSP_OUT_BUF = _param_69FDB_RSP_OUT_BUF;
								// Trace: src/VX_mem_switch.sv:10:15
								localparam ARBITER = _param_69FDB_ARBITER;
								// Trace: src/VX_mem_switch.sv:11:15
								localparam NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? ((NUM_INPUTS + NUM_OUTPUTS) - 1) / NUM_OUTPUTS : ((NUM_OUTPUTS + NUM_INPUTS) - 1) / NUM_INPUTS);
								// Trace: src/VX_mem_switch.sv:12:15
								localparam SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
								// Trace: src/VX_mem_switch.sv:13:15
								localparam LOG_NUM_REQS = $clog2(NUM_REQS);
								// Trace: src/VX_mem_switch.sv:15:5
								wire clk;
								// Trace: src/VX_mem_switch.sv:16:5
								wire reset;
								// Trace: src/VX_mem_switch.sv:17:5
								wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] bus_sel;
								// Trace: src/VX_mem_switch.sv:18:5
								localparam _mbase_bus_in_if = 0;
								// Trace: src/VX_mem_switch.sv:19:5
								localparam _mbase_bus_out_if = 0;
								// Trace: src/VX_mem_switch.sv:21:5
								localparam DATA_WIDTH = 512;
								// Trace: src/VX_mem_switch.sv:22:5
								localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
								localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
								localparam REQ_DATAW = 613;
								// Trace: src/VX_mem_switch.sv:23:5
								localparam RSP_DATAW = 519;
								// Trace: src/VX_mem_switch.sv:24:5
								wire [0:0] req_valid_in;
								// Trace: src/VX_mem_switch.sv:25:5
								wire [612:0] req_data_in;
								// Trace: src/VX_mem_switch.sv:26:5
								wire [0:0] req_ready_in;
								// Trace: src/VX_mem_switch.sv:27:5
								wire [NUM_OUTPUTS - 1:0] req_valid_out;
								// Trace: src/VX_mem_switch.sv:28:5
								wire [(NUM_OUTPUTS * 613) - 1:0] req_data_out;
								// Trace: src/VX_mem_switch.sv:29:5
								wire [NUM_OUTPUTS - 1:0] req_ready_out;
								// Trace: src/VX_mem_switch.sv:30:5
								genvar _gv_i_109;
								for (_gv_i_109 = 0; _gv_i_109 < NUM_INPUTS; _gv_i_109 = _gv_i_109 + 1) begin : g_req_data_in
									localparam i = _gv_i_109;
									// Trace: src/VX_mem_switch.sv:31:9
									assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_bus_in_if].req_valid;
									// Trace: src/VX_mem_switch.sv:32:9
									assign req_data_in[i * 613+:613] = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_bus_in_if].req_data;
									// Trace: src/VX_mem_switch.sv:33:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
								end
								// Trace: src/VX_mem_switch.sv:35:5
								VX_stream_switch #(
									.NUM_INPUTS(NUM_INPUTS),
									.NUM_OUTPUTS(NUM_OUTPUTS),
									.DATAW(REQ_DATAW),
									.OUT_BUF(REQ_OUT_BUF)
								) req_switch(
									.clk(clk),
									.reset(reset),
									.sel_in(bus_sel),
									.valid_in(req_valid_in),
									.data_in(req_data_in),
									.ready_in(req_ready_in),
									.valid_out(req_valid_out),
									.data_out(req_data_out),
									.ready_out(req_ready_out)
								);
								// Trace: src/VX_mem_switch.sv:51:5
								genvar _gv_i_110;
								for (_gv_i_110 = 0; _gv_i_110 < NUM_OUTPUTS; _gv_i_110 = _gv_i_110 + 1) begin : g_req_data_out
									localparam i = _gv_i_110;
									// Trace: src/VX_mem_switch.sv:52:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
									// Trace: src/VX_mem_switch.sv:53:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_data = req_data_out[i * 613+:613];
									// Trace: src/VX_mem_switch.sv:54:9
									assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_ready;
								end
								// Trace: src/VX_mem_switch.sv:56:5
								wire [NUM_OUTPUTS - 1:0] rsp_valid_in;
								// Trace: src/VX_mem_switch.sv:57:5
								wire [(NUM_OUTPUTS * 519) - 1:0] rsp_data_in;
								// Trace: src/VX_mem_switch.sv:58:5
								wire [NUM_OUTPUTS - 1:0] rsp_ready_in;
								// Trace: src/VX_mem_switch.sv:59:5
								wire [0:0] rsp_valid_out;
								// Trace: src/VX_mem_switch.sv:60:5
								wire [518:0] rsp_data_out;
								// Trace: src/VX_mem_switch.sv:61:5
								wire [0:0] rsp_ready_out;
								// Trace: src/VX_mem_switch.sv:62:5
								genvar _gv_i_111;
								for (_gv_i_111 = 0; _gv_i_111 < NUM_OUTPUTS; _gv_i_111 = _gv_i_111 + 1) begin : g_rsp_data_in
									localparam i = _gv_i_111;
									// Trace: src/VX_mem_switch.sv:63:9
									assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_valid;
									// Trace: src/VX_mem_switch.sv:64:9
									assign rsp_data_in[i * 519+:519] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_data;
									// Trace: src/VX_mem_switch.sv:65:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
								end
								// Trace: src/VX_mem_switch.sv:67:5
								VX_stream_arb #(
									.NUM_INPUTS(NUM_OUTPUTS),
									.NUM_OUTPUTS(NUM_INPUTS),
									.DATAW(RSP_DATAW),
									.ARBITER(ARBITER),
									.OUT_BUF(RSP_OUT_BUF)
								) rsp_arb(
									.clk(clk),
									.reset(reset),
									.valid_in(rsp_valid_in),
									.data_in(rsp_data_in),
									.ready_in(rsp_ready_in),
									.valid_out(rsp_valid_out),
									.data_out(rsp_data_out),
									.ready_out(rsp_ready_out),
									.sel_out()
								);
								// Trace: src/VX_mem_switch.sv:84:5
								genvar _gv_i_112;
								for (_gv_i_112 = 0; _gv_i_112 < NUM_INPUTS; _gv_i_112 = _gv_i_112 + 1) begin : g_rsp_data_out
									localparam i = _gv_i_112;
									// Trace: src/VX_mem_switch.sv:85:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
									// Trace: src/VX_mem_switch.sv:86:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 519+:519];
									// Trace: src/VX_mem_switch.sv:87:9
									assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_bus_in_if].rsp_ready;
								end
							end
							assign core_bus_nc_switch.clk = clk;
							assign core_bus_nc_switch.reset = reset;
							assign core_bus_nc_switch.bus_sel = core_req_nc_sel;
							// Trace: src/VX_cache_bypass.sv:58:5
							// expanded interface instance: core_bus_in_nc_if
							localparam _param_C0263_DATA_SIZE = WORD_SIZE;
							localparam _param_C0263_TAG_WIDTH = CORE_TAG_WIDTH;
							genvar _arr_C0263;
							for (_arr_C0263 = 0; _arr_C0263 <= 0; _arr_C0263 = _arr_C0263 + 1) begin : core_bus_in_nc_if
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_C0263_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
								localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
								localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_C0263_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:8:5
								localparam VX_gpu_pkg_UUID_WIDTH = 1;
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:12:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:20:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:24:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire [612:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire [518:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:30:5
								// Trace: src/VX_mem_bus_if.sv:38:5
							end
							// Trace: src/VX_cache_bypass.sv:62:5
							genvar _gv_i_57;
							for (_gv_i_57 = 0; _gv_i_57 < NUM_REQS; _gv_i_57 = _gv_i_57 + 1) begin : g_core_bus_nc_switch_if
								localparam i = _gv_i_57;
								// Trace: src/VX_cache_bypass.sv:63:9
								assign core_bus_in_nc_if[i].req_valid = core_bus_nc_switch_if[0 + i].req_valid;
								// Trace: src/VX_cache_bypass.sv:64:9
								assign core_bus_in_nc_if[i].req_data = core_bus_nc_switch_if[0 + i].req_data;
								// Trace: src/VX_cache_bypass.sv:65:9
								assign core_bus_nc_switch_if[0 + i].req_ready = core_bus_in_nc_if[i].req_ready;
								// Trace: src/VX_cache_bypass.sv:66:9
								assign core_bus_nc_switch_if[0 + i].rsp_valid = core_bus_in_nc_if[i].rsp_valid;
								// Trace: src/VX_cache_bypass.sv:67:9
								assign core_bus_nc_switch_if[0 + i].rsp_data = core_bus_in_nc_if[i].rsp_data;
								// Trace: src/VX_cache_bypass.sv:68:9
								assign core_bus_in_nc_if[i].rsp_ready = core_bus_nc_switch_if[0 + i].rsp_ready;
								if (CACHE_ENABLE) begin : g_cache
									// Trace: src/VX_cache_bypass.sv:70:13
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = core_bus_nc_switch_if[1 + i].req_valid;
									// Trace: src/VX_cache_bypass.sv:71:13
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = core_bus_nc_switch_if[1 + i].req_data;
									// Trace: src/VX_cache_bypass.sv:72:13
									assign core_bus_nc_switch_if[1 + i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_ready;
									// Trace: src/VX_cache_bypass.sv:73:13
									assign core_bus_nc_switch_if[1 + i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_valid;
									// Trace: src/VX_cache_bypass.sv:74:13
									assign core_bus_nc_switch_if[1 + i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_data;
									// Trace: src/VX_cache_bypass.sv:75:13
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = core_bus_nc_switch_if[1 + i].rsp_ready;
								end
								else begin : g_no_cache
									// Trace: src/VX_cache_bypass.sv:77:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = 0;
									// Trace: src/VX_cache_bypass.sv:78:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = 1'sb0;
									// Trace: src/VX_cache_bypass.sv:79:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = 0;
								end
							end
							// Trace: src/VX_cache_bypass.sv:82:5
							// expanded interface instance: core_bus_nc_arb_if
							localparam _param_D50AC_DATA_SIZE = WORD_SIZE;
							localparam _param_D50AC_TAG_WIDTH = MEM_TAG_NC1_WIDTH;
							genvar _arr_D50AC;
							for (_arr_D50AC = 0; _arr_D50AC <= 0; _arr_D50AC = _arr_D50AC + 1) begin : core_bus_nc_arb_if
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_D50AC_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
								localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
								localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_D50AC_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:8:5
								localparam VX_gpu_pkg_UUID_WIDTH = 1;
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:12:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:20:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:24:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire [612:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire [518:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:30:5
								// Trace: src/VX_mem_bus_if.sv:38:5
							end
							// Trace: src/VX_cache_bypass.sv:86:5
							// expanded module instance: core_bus_nc_arb
							localparam _bbase_1376F_bus_in_if = 0;
							localparam _bbase_1376F_bus_out_if = 0;
							localparam _param_1376F_NUM_INPUTS = NUM_REQS;
							localparam _param_1376F_NUM_OUTPUTS = MEM_PORTS;
							localparam _param_1376F_DATA_SIZE = WORD_SIZE;
							localparam _param_1376F_TAG_WIDTH = CORE_TAG_WIDTH;
							localparam _param_1376F_TAG_SEL_IDX = TAG_SEL_IDX;
							localparam _param_1376F_ARBITER = (CACHE_ENABLE ? "P" : "R");
							localparam _param_1376F_REQ_OUT_BUF = 0;
							localparam _param_1376F_RSP_OUT_BUF = 0;
							if (1) begin : core_bus_nc_arb
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_arb.sv:2:15
								localparam NUM_INPUTS = _param_1376F_NUM_INPUTS;
								// Trace: src/VX_mem_arb.sv:3:15
								localparam NUM_OUTPUTS = _param_1376F_NUM_OUTPUTS;
								// Trace: src/VX_mem_arb.sv:4:15
								localparam DATA_SIZE = _param_1376F_DATA_SIZE;
								// Trace: src/VX_mem_arb.sv:5:15
								localparam TAG_WIDTH = _param_1376F_TAG_WIDTH;
								// Trace: src/VX_mem_arb.sv:6:15
								localparam TAG_SEL_IDX = _param_1376F_TAG_SEL_IDX;
								// Trace: src/VX_mem_arb.sv:7:15
								localparam REQ_OUT_BUF = _param_1376F_REQ_OUT_BUF;
								// Trace: src/VX_mem_arb.sv:8:15
								localparam RSP_OUT_BUF = _param_1376F_RSP_OUT_BUF;
								// Trace: src/VX_mem_arb.sv:9:15
								localparam ARBITER = _param_1376F_ARBITER;
								// Trace: src/VX_mem_arb.sv:10:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_arb.sv:11:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_arb.sv:12:15
								localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
								localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
								localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
								// Trace: src/VX_mem_arb.sv:14:5
								wire clk;
								// Trace: src/VX_mem_arb.sv:15:5
								wire reset;
								// Trace: src/VX_mem_arb.sv:16:5
								localparam _mbase_bus_in_if = 0;
								// Trace: src/VX_mem_arb.sv:17:5
								localparam _mbase_bus_out_if = 0;
								// Trace: src/VX_mem_arb.sv:19:5
								localparam DATA_WIDTH = 512;
								// Trace: src/VX_mem_arb.sv:20:5
								localparam LOG_NUM_REQS = 0;
								// Trace: src/VX_mem_arb.sv:21:5
								localparam REQ_DATAW = 613;
								// Trace: src/VX_mem_arb.sv:22:5
								localparam RSP_DATAW = 519;
								// Trace: src/VX_mem_arb.sv:23:5
								localparam SEL_COUNT = NUM_OUTPUTS;
								// Trace: src/VX_mem_arb.sv:24:5
								wire [0:0] req_valid_in;
								// Trace: src/VX_mem_arb.sv:25:5
								wire [612:0] req_data_in;
								// Trace: src/VX_mem_arb.sv:26:5
								wire [0:0] req_ready_in;
								// Trace: src/VX_mem_arb.sv:27:5
								wire [0:0] req_valid_out;
								// Trace: src/VX_mem_arb.sv:28:5
								wire [612:0] req_data_out;
								// Trace: src/VX_mem_arb.sv:29:5
								wire [0:0] req_sel_out;
								// Trace: src/VX_mem_arb.sv:30:5
								wire [0:0] req_ready_out;
								// Trace: src/VX_mem_arb.sv:31:5
								genvar _gv_i_183;
								for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
									localparam i = _gv_i_183;
									// Trace: src/VX_mem_arb.sv:32:9
									assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_valid;
									// Trace: src/VX_mem_arb.sv:33:9
									assign req_data_in[i * 613+:613] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_data;
									// Trace: src/VX_mem_arb.sv:34:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
								end
								// Trace: src/VX_mem_arb.sv:36:5
								VX_stream_arb #(
									.NUM_INPUTS(NUM_INPUTS),
									.NUM_OUTPUTS(NUM_OUTPUTS),
									.DATAW(REQ_DATAW),
									.ARBITER(ARBITER),
									.OUT_BUF(REQ_OUT_BUF)
								) req_arb(
									.clk(clk),
									.reset(reset),
									.valid_in(req_valid_in),
									.ready_in(req_ready_in),
									.data_in(req_data_in),
									.data_out(req_data_out),
									.sel_out(req_sel_out),
									.valid_out(req_valid_out),
									.ready_out(req_ready_out)
								);
								// Trace: src/VX_mem_arb.sv:53:5
								genvar _gv_i_184;
								for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
									localparam i = _gv_i_184;
									// Trace: src/VX_mem_arb.sv:54:9
									wire [6:0] req_tag_out;
									// Trace: src/VX_mem_arb.sv:55:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
									// Trace: src/VX_mem_arb.sv:56:9
									assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[612], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[611-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[585-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[73-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[9-:3], req_tag_out} = req_data_out[i * 613+:613];
									// Trace: src/VX_mem_arb.sv:64:9
									assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_ready;
									if (1) begin : g_req_tag_out
										// Trace: src/VX_mem_arb.sv:76:13
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[6-:7] = req_tag_out;
									end
								end
								// Trace: src/VX_mem_arb.sv:79:5
								wire [0:0] rsp_valid_out;
								// Trace: src/VX_mem_arb.sv:80:5
								wire [518:0] rsp_data_out;
								// Trace: src/VX_mem_arb.sv:81:5
								wire [0:0] rsp_ready_out;
								// Trace: src/VX_mem_arb.sv:82:5
								wire [0:0] rsp_valid_in;
								// Trace: src/VX_mem_arb.sv:83:5
								wire [518:0] rsp_data_in;
								// Trace: src/VX_mem_arb.sv:84:5
								wire [0:0] rsp_ready_in;
								// Trace: src/VX_mem_arb.sv:85:5
								if (1) begin : g_rsp_arb
									genvar _gv_i_186;
									for (_gv_i_186 = 0; _gv_i_186 < NUM_OUTPUTS; _gv_i_186 = _gv_i_186 + 1) begin : g_rsp_data_in
										localparam i = _gv_i_186;
										// Trace: src/VX_mem_arb.sv:120:13
										assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_valid;
										// Trace: src/VX_mem_arb.sv:121:13
										assign rsp_data_in[i * 519+:519] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_data;
										// Trace: src/VX_mem_arb.sv:122:13
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:124:9
									VX_stream_arb #(
										.NUM_INPUTS(NUM_OUTPUTS),
										.NUM_OUTPUTS(NUM_INPUTS),
										.DATAW(RSP_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(RSP_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(rsp_valid_in),
										.ready_in(rsp_ready_in),
										.data_in(rsp_data_in),
										.data_out(rsp_data_out),
										.valid_out(rsp_valid_out),
										.ready_out(rsp_ready_out),
										.sel_out()
									);
								end
								// Trace: src/VX_mem_arb.sv:142:5
								genvar _gv_i_187;
								for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
									localparam i = _gv_i_187;
									// Trace: src/VX_mem_arb.sv:143:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
									// Trace: src/VX_mem_arb.sv:144:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 519+:519];
									// Trace: src/VX_mem_arb.sv:145:9
									assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_ready;
								end
							end
							assign core_bus_nc_arb.clk = clk;
							assign core_bus_nc_arb.reset = reset;
							// Trace: src/VX_cache_bypass.sv:101:5
							// expanded interface instance: mem_bus_out_nc_if
							localparam _param_0061C_DATA_SIZE = LINE_SIZE;
							localparam _param_0061C_TAG_WIDTH = MEM_TAG_NC2_WIDTH;
							genvar _arr_0061C;
							for (_arr_0061C = 0; _arr_0061C <= 0; _arr_0061C = _arr_0061C + 1) begin : mem_bus_out_nc_if
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_0061C_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
								localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
								localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_0061C_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:8:5
								localparam VX_gpu_pkg_UUID_WIDTH = 1;
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:12:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:20:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:24:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire [612:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire [518:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:30:5
								// Trace: src/VX_mem_bus_if.sv:38:5
							end
							// Trace: src/VX_cache_bypass.sv:105:5
							genvar _gv_i_58;
							localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
							localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
							for (_gv_i_58 = 0; _gv_i_58 < MEM_PORTS; _gv_i_58 = _gv_i_58 + 1) begin : g_mem_bus_out_nc
								localparam i = _gv_i_58;
								// Trace: src/VX_cache_bypass.sv:106:9
								wire core_req_nc_arb_rw;
								// Trace: src/VX_cache_bypass.sv:107:9
								wire [63:0] core_req_nc_arb_byteen;
								// Trace: src/VX_cache_bypass.sv:108:9
								wire [25:0] core_req_nc_arb_addr;
								// Trace: src/VX_cache_bypass.sv:109:9
								wire [2:0] core_req_nc_arb_flags;
								// Trace: src/VX_cache_bypass.sv:110:9
								wire [511:0] core_req_nc_arb_data;
								// Trace: src/VX_cache_bypass.sv:111:9
								wire [6:0] core_req_nc_arb_tag;
								// Trace: src/VX_cache_bypass.sv:112:9
								assign {core_req_nc_arb_rw, core_req_nc_arb_addr, core_req_nc_arb_data, core_req_nc_arb_byteen, core_req_nc_arb_flags, core_req_nc_arb_tag} = core_bus_nc_arb_if[i].req_data;
								// Trace: src/VX_cache_bypass.sv:120:9
								wire [25:0] core_req_nc_arb_addr_w;
								// Trace: src/VX_cache_bypass.sv:121:9
								wire [63:0] core_req_nc_arb_byteen_w;
								// Trace: src/VX_cache_bypass.sv:122:9
								wire [511:0] core_req_nc_arb_data_w;
								// Trace: src/VX_cache_bypass.sv:123:9
								wire [511:0] core_rsp_nc_arb_data_w;
								// Trace: src/VX_cache_bypass.sv:124:9
								wire [6:0] core_req_nc_arb_tag_w;
								// Trace: src/VX_cache_bypass.sv:125:9
								wire [6:0] core_rsp_nc_arb_tag_w;
								if (1) begin : g_single_word_line
									// Trace: src/VX_cache_bypass.sv:156:13
									assign core_req_nc_arb_addr_w = core_req_nc_arb_addr;
									// Trace: src/VX_cache_bypass.sv:157:13
									assign core_req_nc_arb_byteen_w = core_req_nc_arb_byteen;
									// Trace: src/VX_cache_bypass.sv:158:13
									assign core_req_nc_arb_data_w = core_req_nc_arb_data;
									// Trace: src/VX_cache_bypass.sv:159:13
									assign core_req_nc_arb_tag_w = core_req_nc_arb_tag;
									// Trace: src/VX_cache_bypass.sv:160:13
									assign core_rsp_nc_arb_data_w = mem_bus_out_nc_if[i].rsp_data[518-:512];
									// Trace: src/VX_cache_bypass.sv:161:13
									assign core_rsp_nc_arb_tag_w = sv2v_cast_7(mem_bus_out_nc_if[i].rsp_data[6-:7]);
								end
								// Trace: src/VX_cache_bypass.sv:163:9
								assign mem_bus_out_nc_if[i].req_valid = core_bus_nc_arb_if[i].req_valid;
								// Trace: src/VX_cache_bypass.sv:164:9
								assign mem_bus_out_nc_if[i].req_data = {core_req_nc_arb_rw, core_req_nc_arb_addr_w, core_req_nc_arb_data_w, core_req_nc_arb_byteen_w, core_req_nc_arb_flags, core_req_nc_arb_tag_w};
								// Trace: src/VX_cache_bypass.sv:172:9
								assign core_bus_nc_arb_if[i].req_ready = mem_bus_out_nc_if[i].req_ready;
								// Trace: src/VX_cache_bypass.sv:173:9
								assign core_bus_nc_arb_if[i].rsp_valid = mem_bus_out_nc_if[i].rsp_valid;
								// Trace: src/VX_cache_bypass.sv:174:9
								assign core_bus_nc_arb_if[i].rsp_data = {core_rsp_nc_arb_data_w, core_rsp_nc_arb_tag_w};
								// Trace: src/VX_cache_bypass.sv:178:9
								assign mem_bus_out_nc_if[i].rsp_ready = core_bus_nc_arb_if[i].rsp_ready;
							end
							// Trace: src/VX_cache_bypass.sv:180:5
							// expanded interface instance: mem_bus_out_src_if
							localparam _param_913F6_DATA_SIZE = LINE_SIZE;
							localparam _param_913F6_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
							genvar _arr_913F6;
							for (_arr_913F6 = 0; _arr_913F6 <= (((CACHE_ENABLE ? 2 : 1) * MEM_PORTS) - 1); _arr_913F6 = _arr_913F6 + 1) begin : mem_bus_out_src_if
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_913F6_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
								localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
								localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_913F6_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:8:5
								localparam VX_gpu_pkg_UUID_WIDTH = 1;
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:12:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:20:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:24:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire [612:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire [518:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:30:5
								// Trace: src/VX_mem_bus_if.sv:38:5
							end
							// Trace: src/VX_cache_bypass.sv:184:5
							genvar _gv_i_59;
							for (_gv_i_59 = 0; _gv_i_59 < MEM_PORTS; _gv_i_59 = _gv_i_59 + 1) begin : g_mem_bus_out_src
								localparam i = _gv_i_59;
								// Trace: src/VX_cache_bypass.sv:186:5
								assign mem_bus_out_src_if[0 + i].req_valid = mem_bus_out_nc_if[i].req_valid;
								// Trace: src/VX_cache_bypass.sv:187:5
								assign mem_bus_out_src_if[0 + i].req_data[612] = mem_bus_out_nc_if[i].req_data[612];
								// Trace: src/VX_cache_bypass.sv:188:5
								assign mem_bus_out_src_if[0 + i].req_data[611-:26] = mem_bus_out_nc_if[i].req_data[611-:26];
								// Trace: src/VX_cache_bypass.sv:189:5
								assign mem_bus_out_src_if[0 + i].req_data[585-:512] = mem_bus_out_nc_if[i].req_data[585-:512];
								// Trace: src/VX_cache_bypass.sv:190:5
								assign mem_bus_out_src_if[0 + i].req_data[73-:64] = mem_bus_out_nc_if[i].req_data[73-:64];
								// Trace: src/VX_cache_bypass.sv:191:5
								assign mem_bus_out_src_if[0 + i].req_data[9-:3] = mem_bus_out_nc_if[i].req_data[9-:3];
								if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk1
									if (1) begin : genblk1
										if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
											// Trace: src/VX_cache_bypass.sv:195:17
											assign mem_bus_out_src_if[0 + i].req_data[6-:7] = {mem_bus_out_nc_if[i].req_data[6-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_NC2_WIDTH {1'b0}}, mem_bus_out_nc_if[i].req_data[5-:6]};
										end
										else begin : genblk1
											// Trace: src/VX_cache_bypass.sv:197:17
											assign mem_bus_out_src_if[0 + i].req_data[6-:7] = {mem_bus_out_nc_if[i].req_data[6-:1], mem_bus_out_nc_if[i].req_data[(MEM_TAG_OUT_WIDTH - VX_gpu_pkg_UUID_WIDTH) - 1:0]};
										end
									end
								end
								else begin : genblk1
									// Trace: src/VX_cache_bypass.sv:207:9
									assign mem_bus_out_src_if[0 + i].req_data[6-:7] = mem_bus_out_nc_if[i].req_data[6-:7];
								end
								// Trace: src/VX_cache_bypass.sv:209:5
								assign mem_bus_out_nc_if[i].req_ready = mem_bus_out_src_if[0 + i].req_ready;
								// Trace: src/VX_cache_bypass.sv:210:5
								assign mem_bus_out_nc_if[i].rsp_valid = mem_bus_out_src_if[0 + i].rsp_valid;
								// Trace: src/VX_cache_bypass.sv:211:5
								assign mem_bus_out_nc_if[i].rsp_data[518-:512] = mem_bus_out_src_if[0 + i].rsp_data[518-:512];
								if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk2
									if (1) begin : genblk1
										if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
											// Trace: src/VX_cache_bypass.sv:215:17
											assign mem_bus_out_nc_if[i].rsp_data[6-:7] = {mem_bus_out_src_if[0 + i].rsp_data[6-:1], mem_bus_out_src_if[0 + i].rsp_data[5:0]};
										end
										else begin : genblk1
											// Trace: src/VX_cache_bypass.sv:217:17
											assign mem_bus_out_nc_if[i].rsp_data[6-:7] = {mem_bus_out_src_if[0 + i].rsp_data[6-:1], {MEM_TAG_NC2_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[0 + i].rsp_data[5-:6]};
										end
									end
								end
								else begin : genblk2
									// Trace: src/VX_cache_bypass.sv:227:9
									assign mem_bus_out_nc_if[i].rsp_data[6-:7] = mem_bus_out_src_if[0 + i].rsp_data[6-:7];
								end
								// Trace: src/VX_cache_bypass.sv:229:5
								assign mem_bus_out_src_if[0 + i].rsp_ready = mem_bus_out_nc_if[i].rsp_ready;
								if (CACHE_ENABLE) begin : g_cache
									// Trace: src/VX_cache_bypass.sv:233:5
									assign mem_bus_out_src_if[1 + i].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_valid;
									// Trace: src/VX_cache_bypass.sv:234:5
									assign mem_bus_out_src_if[1 + i].req_data[612] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[610];
									// Trace: src/VX_cache_bypass.sv:235:5
									assign mem_bus_out_src_if[1 + i].req_data[611-:26] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[609-:26];
									// Trace: src/VX_cache_bypass.sv:236:5
									assign mem_bus_out_src_if[1 + i].req_data[585-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[583-:512];
									// Trace: src/VX_cache_bypass.sv:237:5
									assign mem_bus_out_src_if[1 + i].req_data[73-:64] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[71-:64];
									// Trace: src/VX_cache_bypass.sv:238:5
									assign mem_bus_out_src_if[1 + i].req_data[9-:3] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[7-:3];
									if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk1
										if (1) begin : genblk1
											if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
												// Trace: src/VX_cache_bypass.sv:242:17
												assign mem_bus_out_src_if[1 + i].req_data[6-:7] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_IN_WIDTH {1'b0}}, Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[3-:4]};
											end
											else begin : genblk1
												// Trace: src/VX_cache_bypass.sv:244:17
												assign mem_bus_out_src_if[1 + i].req_data[6-:7] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[(MEM_TAG_OUT_WIDTH - VX_gpu_pkg_UUID_WIDTH) - 1:0]};
											end
										end
									end
									else begin : genblk1
										// Trace: src/VX_cache_bypass.sv:254:9
										assign mem_bus_out_src_if[1 + i].req_data[6-:7] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:5];
									end
									// Trace: src/VX_cache_bypass.sv:256:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = mem_bus_out_src_if[1 + i].req_ready;
									// Trace: src/VX_cache_bypass.sv:257:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = mem_bus_out_src_if[1 + i].rsp_valid;
									// Trace: src/VX_cache_bypass.sv:258:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[516-:512] = mem_bus_out_src_if[1 + i].rsp_data[518-:512];
									if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk2
										if (1) begin : genblk1
											if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
												// Trace: src/VX_cache_bypass.sv:262:17
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[6-:1], mem_bus_out_src_if[1 + i].rsp_data[3:0]};
											end
											else begin : genblk1
												// Trace: src/VX_cache_bypass.sv:264:17
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[6-:1], {MEM_TAG_IN_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[1 + i].rsp_data[5-:6]};
											end
										end
									end
									else begin : genblk2
										// Trace: src/VX_cache_bypass.sv:274:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = mem_bus_out_src_if[1 + i].rsp_data[6-:7];
									end
									// Trace: src/VX_cache_bypass.sv:276:5
									assign mem_bus_out_src_if[1 + i].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_ready;
								end
								else begin : g_no_cache
									// Trace: src/VX_cache_bypass.sv:279:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = 0;
									// Trace: src/VX_cache_bypass.sv:280:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = 0;
									// Trace: src/VX_cache_bypass.sv:281:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data = 1'sb0;
								end
							end
							// Trace: src/VX_cache_bypass.sv:284:5
							// expanded module instance: mem_bus_out_arb
							localparam _bbase_B06D0_bus_in_if = 0;
							localparam _bbase_B06D0_bus_out_if = 0;
							localparam _param_B06D0_NUM_INPUTS = (CACHE_ENABLE ? 2 : 1) * MEM_PORTS;
							localparam _param_B06D0_NUM_OUTPUTS = MEM_PORTS;
							localparam _param_B06D0_DATA_SIZE = LINE_SIZE;
							localparam _param_B06D0_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
							localparam _param_B06D0_ARBITER = "R";
							localparam _param_B06D0_REQ_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
							localparam _param_B06D0_RSP_OUT_BUF = 0;
							if (1) begin : mem_bus_out_arb
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_arb.sv:2:15
								localparam NUM_INPUTS = _param_B06D0_NUM_INPUTS;
								// Trace: src/VX_mem_arb.sv:3:15
								localparam NUM_OUTPUTS = _param_B06D0_NUM_OUTPUTS;
								// Trace: src/VX_mem_arb.sv:4:15
								localparam DATA_SIZE = _param_B06D0_DATA_SIZE;
								// Trace: src/VX_mem_arb.sv:5:15
								localparam TAG_WIDTH = _param_B06D0_TAG_WIDTH;
								// Trace: src/VX_mem_arb.sv:6:15
								localparam TAG_SEL_IDX = 0;
								// Trace: src/VX_mem_arb.sv:7:15
								localparam REQ_OUT_BUF = _param_B06D0_REQ_OUT_BUF;
								// Trace: src/VX_mem_arb.sv:8:15
								localparam RSP_OUT_BUF = _param_B06D0_RSP_OUT_BUF;
								// Trace: src/VX_mem_arb.sv:9:15
								localparam ARBITER = _param_B06D0_ARBITER;
								// Trace: src/VX_mem_arb.sv:10:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_arb.sv:11:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_arb.sv:12:15
								localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
								localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
								localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
								// Trace: src/VX_mem_arb.sv:14:5
								wire clk;
								// Trace: src/VX_mem_arb.sv:15:5
								wire reset;
								// Trace: src/VX_mem_arb.sv:16:5
								localparam _mbase_bus_in_if = 0;
								// Trace: src/VX_mem_arb.sv:17:5
								localparam _mbase_bus_out_if = 0;
								// Trace: src/VX_mem_arb.sv:19:5
								localparam DATA_WIDTH = 512;
								// Trace: src/VX_mem_arb.sv:20:5
								localparam LOG_NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? $clog2((NUM_INPUTS + 0) / 1) : 0);
								// Trace: src/VX_mem_arb.sv:21:5
								localparam REQ_DATAW = 606 + TAG_WIDTH;
								// Trace: src/VX_mem_arb.sv:22:5
								localparam RSP_DATAW = DATA_WIDTH + TAG_WIDTH;
								// Trace: src/VX_mem_arb.sv:23:5
								localparam SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
								// Trace: src/VX_mem_arb.sv:24:5
								wire [NUM_INPUTS - 1:0] req_valid_in;
								// Trace: src/VX_mem_arb.sv:25:5
								wire [(NUM_INPUTS * REQ_DATAW) - 1:0] req_data_in;
								// Trace: src/VX_mem_arb.sv:26:5
								wire [NUM_INPUTS - 1:0] req_ready_in;
								// Trace: src/VX_mem_arb.sv:27:5
								wire [0:0] req_valid_out;
								// Trace: src/VX_mem_arb.sv:28:5
								wire [REQ_DATAW - 1:0] req_data_out;
								// Trace: src/VX_mem_arb.sv:29:5
								wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] req_sel_out;
								// Trace: src/VX_mem_arb.sv:30:5
								wire [0:0] req_ready_out;
								// Trace: src/VX_mem_arb.sv:31:5
								genvar _gv_i_183;
								for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
									localparam i = _gv_i_183;
									// Trace: src/VX_mem_arb.sv:32:9
									assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_valid;
									// Trace: src/VX_mem_arb.sv:33:9
									assign req_data_in[i * 613+:613] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_data;
									// Trace: src/VX_mem_arb.sv:34:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
								end
								// Trace: src/VX_mem_arb.sv:36:5
								VX_stream_arb #(
									.NUM_INPUTS(NUM_INPUTS),
									.NUM_OUTPUTS(NUM_OUTPUTS),
									.DATAW(REQ_DATAW),
									.ARBITER(ARBITER),
									.OUT_BUF(REQ_OUT_BUF)
								) req_arb(
									.clk(clk),
									.reset(reset),
									.valid_in(req_valid_in),
									.ready_in(req_ready_in),
									.data_in(req_data_in),
									.data_out(req_data_out),
									.sel_out(req_sel_out),
									.valid_out(req_valid_out),
									.ready_out(req_ready_out)
								);
								// Trace: src/VX_mem_arb.sv:53:5
								genvar _gv_i_184;
								for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
									localparam i = _gv_i_184;
									// Trace: src/VX_mem_arb.sv:54:9
									wire [TAG_WIDTH - 1:0] req_tag_out;
									// Trace: src/VX_mem_arb.sv:55:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
									// Trace: src/VX_mem_arb.sv:56:9
									assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[612], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[611-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[585-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[73-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[9-:3], req_tag_out} = req_data_out[i * 613+:613];
									// Trace: src/VX_mem_arb.sv:64:9
									assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
									if (NUM_INPUTS > NUM_OUTPUTS) begin : g_req_tag_sel_out
										// Trace: src/VX_mem_arb.sv:66:13
										VX_bits_insert #(
											.N(TAG_WIDTH),
											.S(LOG_NUM_REQS),
											.POS(TAG_SEL_IDX)
										) bits_insert(
											.data_in(req_tag_out),
											.ins_in(req_sel_out[i * 1+:1]),
											.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[6-:7])
										);
									end
									else begin : g_req_tag_out
										// Trace: src/VX_mem_arb.sv:76:13
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[6-:7] = req_tag_out;
									end
								end
								// Trace: src/VX_mem_arb.sv:79:5
								wire [NUM_INPUTS - 1:0] rsp_valid_out;
								// Trace: src/VX_mem_arb.sv:80:5
								wire [(NUM_INPUTS * RSP_DATAW) - 1:0] rsp_data_out;
								// Trace: src/VX_mem_arb.sv:81:5
								wire [NUM_INPUTS - 1:0] rsp_ready_out;
								// Trace: src/VX_mem_arb.sv:82:5
								wire [0:0] rsp_valid_in;
								// Trace: src/VX_mem_arb.sv:83:5
								wire [RSP_DATAW - 1:0] rsp_data_in;
								// Trace: src/VX_mem_arb.sv:84:5
								wire [0:0] rsp_ready_in;
								// Trace: src/VX_mem_arb.sv:85:5
								if (NUM_INPUTS > NUM_OUTPUTS) begin : g_rsp_select
									// Trace: src/VX_mem_arb.sv:86:9
									wire [LOG_NUM_REQS - 1:0] rsp_sel_in;
									genvar _gv_i_185;
									for (_gv_i_185 = 0; _gv_i_185 < NUM_OUTPUTS; _gv_i_185 = _gv_i_185 + 1) begin : g_rsp_data_in
										localparam i = _gv_i_185;
										// Trace: src/VX_mem_arb.sv:88:13
										wire [TAG_WIDTH - 1:0] rsp_tag_out;
										// Trace: src/VX_mem_arb.sv:89:13
										VX_bits_remove #(
											.N(TAG_WIDTH + LOG_NUM_REQS),
											.S(LOG_NUM_REQS),
											.POS(TAG_SEL_IDX)
										) bits_remove(
											.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[6-:7]),
											.sel_out(rsp_sel_in[0+:0]),
											.data_out(rsp_tag_out)
										);
										// Trace: src/VX_mem_arb.sv:98:13
										assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
										// Trace: src/VX_mem_arb.sv:99:13
										assign rsp_data_in[i * 519+:519] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[518-:512], rsp_tag_out};
										// Trace: src/VX_mem_arb.sv:100:13
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:102:9
									VX_stream_switch #(
										.NUM_INPUTS(NUM_OUTPUTS),
										.NUM_OUTPUTS(NUM_INPUTS),
										.DATAW(RSP_DATAW),
										.OUT_BUF(RSP_OUT_BUF)
									) rsp_switch(
										.clk(clk),
										.reset(reset),
										.sel_in(rsp_sel_in),
										.valid_in(rsp_valid_in),
										.ready_in(rsp_ready_in),
										.data_in(rsp_data_in),
										.data_out(rsp_data_out),
										.valid_out(rsp_valid_out),
										.ready_out(rsp_ready_out)
									);
								end
								else begin : g_rsp_arb
									genvar _gv_i_186;
									for (_gv_i_186 = 0; _gv_i_186 < NUM_OUTPUTS; _gv_i_186 = _gv_i_186 + 1) begin : g_rsp_data_in
										localparam i = _gv_i_186;
										// Trace: src/VX_mem_arb.sv:120:13
										assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
										// Trace: src/VX_mem_arb.sv:121:13
										assign rsp_data_in[i * 519+:519] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
										// Trace: src/VX_mem_arb.sv:122:13
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:124:9
									VX_stream_arb #(
										.NUM_INPUTS(NUM_OUTPUTS),
										.NUM_OUTPUTS(NUM_INPUTS),
										.DATAW(RSP_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(RSP_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(rsp_valid_in),
										.ready_in(rsp_ready_in),
										.data_in(rsp_data_in),
										.data_out(rsp_data_out),
										.valid_out(rsp_valid_out),
										.ready_out(rsp_ready_out),
										.sel_out()
									);
								end
								// Trace: src/VX_mem_arb.sv:142:5
								genvar _gv_i_187;
								for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
									localparam i = _gv_i_187;
									// Trace: src/VX_mem_arb.sv:143:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
									// Trace: src/VX_mem_arb.sv:144:9
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 519+:519];
									// Trace: src/VX_mem_arb.sv:145:9
									assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.l2cache.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_ready;
								end
							end
							assign mem_bus_out_arb.clk = clk;
							assign mem_bus_out_arb.reset = reset;
						end
						assign cache_bypass.clk = clk;
						assign cache_bypass.reset = reset;
					end
					else begin : g_no_bypass
						genvar _gv_i_38;
						for (_gv_i_38 = 0; _gv_i_38 < NUM_REQS; _gv_i_38 = _gv_i_38 + 1) begin : g_core_bus_cache_if
							localparam i = _gv_i_38;
							// Trace: src/VX_cache_wrap.sv:73:5
							assign core_bus_cache_if[i].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_if].req_valid;
							// Trace: src/VX_cache_wrap.sv:74:5
							assign core_bus_cache_if[i].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_if].req_data;
							// Trace: src/VX_cache_wrap.sv:75:5
							assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_if].req_ready = core_bus_cache_if[i].req_ready;
							// Trace: src/VX_cache_wrap.sv:76:5
							assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_if].rsp_valid = core_bus_cache_if[i].rsp_valid;
							// Trace: src/VX_cache_wrap.sv:77:5
							assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_if].rsp_data = core_bus_cache_if[i].rsp_data;
							// Trace: src/VX_cache_wrap.sv:78:5
							assign core_bus_cache_if[i].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_core_bus_if].rsp_ready;
						end
						genvar _gv_i_39;
						for (_gv_i_39 = 0; _gv_i_39 < MEM_PORTS; _gv_i_39 = _gv_i_39 + 1) begin : g_mem_bus_tmp_if
							localparam i = _gv_i_39;
							// Trace: src/VX_cache_wrap.sv:81:5
							assign mem_bus_tmp_if[i].req_valid = mem_bus_cache_if[i].req_valid;
							// Trace: src/VX_cache_wrap.sv:82:5
							assign mem_bus_tmp_if[i].req_data = mem_bus_cache_if[i].req_data;
							// Trace: src/VX_cache_wrap.sv:83:5
							assign mem_bus_cache_if[i].req_ready = mem_bus_tmp_if[i].req_ready;
							// Trace: src/VX_cache_wrap.sv:84:5
							assign mem_bus_cache_if[i].rsp_valid = mem_bus_tmp_if[i].rsp_valid;
							// Trace: src/VX_cache_wrap.sv:85:5
							assign mem_bus_cache_if[i].rsp_data = mem_bus_tmp_if[i].rsp_data;
							// Trace: src/VX_cache_wrap.sv:86:5
							assign mem_bus_tmp_if[i].rsp_ready = mem_bus_cache_if[i].rsp_ready;
						end
					end
					// Trace: src/VX_cache_wrap.sv:89:5
					genvar _gv_i_40;
					for (_gv_i_40 = 0; _gv_i_40 < MEM_PORTS; _gv_i_40 = _gv_i_40 + 1) begin : g_mem_bus_if
						localparam i = _gv_i_40;
						if (WRITE_ENABLE) begin : g_we
							// Trace: src/VX_cache_wrap.sv:91:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
							// Trace: src/VX_cache_wrap.sv:92:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[i].req_data;
							// Trace: src/VX_cache_wrap.sv:93:5
							assign mem_bus_tmp_if[i].req_ready = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
							// Trace: src/VX_cache_wrap.sv:94:5
							assign mem_bus_tmp_if[i].rsp_valid = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
							// Trace: src/VX_cache_wrap.sv:95:5
							assign mem_bus_tmp_if[i].rsp_data = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
							// Trace: src/VX_cache_wrap.sv:96:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
						end
						else begin : g_ro
							// Trace: src/VX_cache_wrap.sv:98:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
							// Trace: src/VX_cache_wrap.sv:99:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data[612] = 0;
							// Trace: src/VX_cache_wrap.sv:100:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data[611-:26] = mem_bus_tmp_if[i].req_data[611-:26];
							// Trace: src/VX_cache_wrap.sv:101:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data[585-:512] = 1'sb0;
							// Trace: src/VX_cache_wrap.sv:102:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data[73-:64] = 1'sb1;
							// Trace: src/VX_cache_wrap.sv:103:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data[9-:3] = mem_bus_tmp_if[i].req_data[9-:3];
							// Trace: src/VX_cache_wrap.sv:104:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_data[6-:7] = mem_bus_tmp_if[i].req_data[6-:7];
							// Trace: src/VX_cache_wrap.sv:105:5
							assign mem_bus_tmp_if[i].req_ready = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
							// Trace: src/VX_cache_wrap.sv:106:5
							assign mem_bus_tmp_if[i].rsp_valid = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
							// Trace: src/VX_cache_wrap.sv:107:5
							assign mem_bus_tmp_if[i].rsp_data[518-:512] = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[518-:512];
							// Trace: src/VX_cache_wrap.sv:108:5
							assign mem_bus_tmp_if[i].rsp_data[6-:7] = Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[6-:7];
							// Trace: src/VX_cache_wrap.sv:109:5
							assign Vortex.per_cluster_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
						end
					end
					// Trace: src/VX_cache_wrap.sv:112:5
					if (1) begin : g_passthru
						genvar _gv_i_41;
						for (_gv_i_41 = 0; _gv_i_41 < NUM_REQS; _gv_i_41 = _gv_i_41 + 1) begin : g_core_bus_cache_if
							localparam i = _gv_i_41;
							// Trace: src/VX_cache_wrap.sv:141:5
							assign core_bus_cache_if[i].req_ready = 0;
							// Trace: src/VX_cache_wrap.sv:142:5
							assign core_bus_cache_if[i].rsp_valid = 0;
							// Trace: src/VX_cache_wrap.sv:143:5
							assign core_bus_cache_if[i].rsp_data = 1'sb0;
						end
						genvar _gv_i_42;
						for (_gv_i_42 = 0; _gv_i_42 < MEM_PORTS; _gv_i_42 = _gv_i_42 + 1) begin : g_mem_bus_cache_if
							localparam i = _gv_i_42;
							// Trace: src/VX_cache_wrap.sv:146:5
							assign mem_bus_cache_if[i].req_valid = 0;
							// Trace: src/VX_cache_wrap.sv:147:5
							assign mem_bus_cache_if[i].req_data = 1'sb0;
							// Trace: src/VX_cache_wrap.sv:148:5
							assign mem_bus_cache_if[i].rsp_ready = 0;
						end
					end
				end
				assign l2cache.clk = clk;
				assign l2cache.reset = l2_reset;
				// Trace: src/VX_cluster.sv:49:5
				wire [0:0] per_socket_busy;
				// Trace: src/VX_cluster.sv:50:5
				genvar _gv_socket_id_1;
				localparam VX_gpu_pkg_VX_DCR_ADDR_WIDTH = 12;
				localparam VX_gpu_pkg_VX_DCR_DATA_WIDTH = 32;
				for (_gv_socket_id_1 = 0; _gv_socket_id_1 < VX_gpu_pkg_NUM_SOCKETS; _gv_socket_id_1 = _gv_socket_id_1 + 1) begin : g_sockets
					localparam socket_id = _gv_socket_id_1;
					// Trace: src/VX_cluster.sv:51:5
					wire [0:0] socket_reset;
					// Trace: src/VX_cluster.sv:52:5
					VX_reset_relay #(
						.N(1),
						.MAX_FANOUT(0)
					) __socket_reset(
						.clk(clk),
						.reset(reset),
						.reset_o(socket_reset)
					);
					// Trace: src/VX_cluster.sv:57:9
					// expanded interface instance: socket_dcr_bus_if
					if (1) begin : socket_dcr_bus_if
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_dcr_bus_if.sv:2:5
						wire write_valid;
						// Trace: src/VX_dcr_bus_if.sv:3:5
						localparam VX_gpu_pkg_VX_DCR_ADDR_WIDTH = 12;
						wire [11:0] write_addr;
						// Trace: src/VX_dcr_bus_if.sv:4:5
						localparam VX_gpu_pkg_VX_DCR_DATA_WIDTH = 32;
						wire [31:0] write_data;
						// Trace: src/VX_dcr_bus_if.sv:5:5
						// Trace: src/VX_dcr_bus_if.sv:10:5
					end
					// Trace: src/VX_cluster.sv:58:9
					wire is_base_dcr_addr = (Vortex.g_clusters[_gv_cluster_id_1].cluster_dcr_bus_if.write_addr >= 12'h001) && (Vortex.g_clusters[_gv_cluster_id_1].cluster_dcr_bus_if.write_addr < 12'h006);
					if (1) begin : genblk1
						// Trace: src/VX_cluster.sv:72:9
						assign {socket_dcr_bus_if.write_valid, socket_dcr_bus_if.write_addr, socket_dcr_bus_if.write_data} = {Vortex.g_clusters[_gv_cluster_id_1].cluster_dcr_bus_if.write_valid && is_base_dcr_addr, Vortex.g_clusters[_gv_cluster_id_1].cluster_dcr_bus_if.write_addr, Vortex.g_clusters[_gv_cluster_id_1].cluster_dcr_bus_if.write_data};
					end
					// Trace: src/VX_cluster.sv:75:9
					// expanded module instance: socket
					localparam _bbase_66BD2_mem_bus_if = socket_id * VX_gpu_pkg_DCACHE_NUM_REQS;
					localparam _param_66BD2_SOCKET_ID = (CLUSTER_ID * VX_gpu_pkg_NUM_SOCKETS) + socket_id;
					localparam _param_66BD2_INSTANCE_ID = "";
					if (1) begin : socket
						// removed import VX_gpu_pkg::*;
						// Trace: src/VX_socket.sv:2:15
						localparam SOCKET_ID = _param_66BD2_SOCKET_ID;
						// Trace: src/VX_socket.sv:3:15
						localparam INSTANCE_ID = _param_66BD2_INSTANCE_ID;
						// Trace: src/VX_socket.sv:5:5
						wire clk;
						// Trace: src/VX_socket.sv:6:5
						wire reset;
						// Trace: src/VX_socket.sv:7:5
						// removed modport instance dcr_bus_if
						// Trace: src/VX_socket.sv:8:5
						localparam VX_gpu_pkg_DCACHE_WORD_SIZE = 16;
						localparam VX_gpu_pkg_XLENB = 4;
						localparam VX_gpu_pkg_LSU_WORD_SIZE = VX_gpu_pkg_XLENB;
						localparam VX_gpu_pkg_DCACHE_CHANNELS = 1;
						localparam VX_gpu_pkg_DCACHE_NUM_REQS = 1;
						localparam _mbase_mem_bus_if = _bbase_66BD2_mem_bus_if;
						// Trace: src/VX_socket.sv:9:5
						wire busy;
						// Trace: src/VX_socket.sv:11:5
						localparam VX_gpu_pkg_NW_BITS = 2;
						localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
						localparam VX_gpu_pkg_ICACHE_TAG_ID_BITS = VX_gpu_pkg_NW_WIDTH;
						localparam VX_gpu_pkg_UUID_WIDTH = 1;
						localparam VX_gpu_pkg_ICACHE_TAG_WIDTH = 3;
						localparam VX_gpu_pkg_ICACHE_WORD_SIZE = 4;
						// expanded interface instance: per_core_icache_bus_if
						localparam _param_FD2E2_DATA_SIZE = VX_gpu_pkg_ICACHE_WORD_SIZE;
						localparam _param_FD2E2_TAG_WIDTH = VX_gpu_pkg_ICACHE_TAG_WIDTH;
						genvar _arr_FD2E2;
						for (_arr_FD2E2 = 0; _arr_FD2E2 <= 0; _arr_FD2E2 = _arr_FD2E2 + 1) begin : per_core_icache_bus_if
							// removed import VX_gpu_pkg::*;
							// Trace: src/VX_mem_bus_if.sv:2:15
							localparam DATA_SIZE = _param_FD2E2_DATA_SIZE;
							// Trace: src/VX_mem_bus_if.sv:3:15
							localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
							localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
							localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
							// Trace: src/VX_mem_bus_if.sv:4:15
							localparam TAG_WIDTH = _param_FD2E2_TAG_WIDTH;
							// Trace: src/VX_mem_bus_if.sv:5:15
							localparam MEM_ADDR_WIDTH = 32;
							// Trace: src/VX_mem_bus_if.sv:6:15
							localparam ADDR_WIDTH = 30;
							// Trace: src/VX_mem_bus_if.sv:8:5
							localparam VX_gpu_pkg_UUID_WIDTH = 1;
							// removed localparam type tag_t
							// Trace: src/VX_mem_bus_if.sv:12:5
							// removed localparam type req_data_t
							// Trace: src/VX_mem_bus_if.sv:20:5
							// removed localparam type rsp_data_t
							// Trace: src/VX_mem_bus_if.sv:24:5
							wire req_valid;
							// Trace: src/VX_mem_bus_if.sv:25:5
							wire [72:0] req_data;
							// Trace: src/VX_mem_bus_if.sv:26:5
							wire req_ready;
							// Trace: src/VX_mem_bus_if.sv:27:5
							wire rsp_valid;
							// Trace: src/VX_mem_bus_if.sv:28:5
							wire [34:0] rsp_data;
							// Trace: src/VX_mem_bus_if.sv:29:5
							wire rsp_ready;
							// Trace: src/VX_mem_bus_if.sv:30:5
							// Trace: src/VX_mem_bus_if.sv:38:5
						end
						// Trace: src/VX_socket.sv:15:5
						localparam VX_gpu_pkg_ICACHE_LINE_SIZE = 64;
						localparam VX_gpu_pkg_ICACHE_MEM_TAG_WIDTH = 5;
						// expanded interface instance: icache_mem_bus_if
						localparam _param_063FD_DATA_SIZE = VX_gpu_pkg_ICACHE_LINE_SIZE;
						localparam _param_063FD_TAG_WIDTH = VX_gpu_pkg_ICACHE_MEM_TAG_WIDTH;
						genvar _arr_063FD;
						for (_arr_063FD = 0; _arr_063FD <= 0; _arr_063FD = _arr_063FD + 1) begin : icache_mem_bus_if
							// removed import VX_gpu_pkg::*;
							// Trace: src/VX_mem_bus_if.sv:2:15
							localparam DATA_SIZE = _param_063FD_DATA_SIZE;
							// Trace: src/VX_mem_bus_if.sv:3:15
							localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
							localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
							localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
							// Trace: src/VX_mem_bus_if.sv:4:15
							localparam TAG_WIDTH = _param_063FD_TAG_WIDTH;
							// Trace: src/VX_mem_bus_if.sv:5:15
							localparam MEM_ADDR_WIDTH = 32;
							// Trace: src/VX_mem_bus_if.sv:6:15
							localparam ADDR_WIDTH = 26;
							// Trace: src/VX_mem_bus_if.sv:8:5
							localparam VX_gpu_pkg_UUID_WIDTH = 1;
							// removed localparam type tag_t
							// Trace: src/VX_mem_bus_if.sv:12:5
							// removed localparam type req_data_t
							// Trace: src/VX_mem_bus_if.sv:20:5
							// removed localparam type rsp_data_t
							// Trace: src/VX_mem_bus_if.sv:24:5
							wire req_valid;
							// Trace: src/VX_mem_bus_if.sv:25:5
							wire [610:0] req_data;
							// Trace: src/VX_mem_bus_if.sv:26:5
							wire req_ready;
							// Trace: src/VX_mem_bus_if.sv:27:5
							wire rsp_valid;
							// Trace: src/VX_mem_bus_if.sv:28:5
							wire [516:0] rsp_data;
							// Trace: src/VX_mem_bus_if.sv:29:5
							wire rsp_ready;
							// Trace: src/VX_mem_bus_if.sv:30:5
							// Trace: src/VX_mem_bus_if.sv:38:5
						end
						// Trace: src/VX_socket.sv:19:5
						wire [0:0] icache_reset;
						// Trace: src/VX_socket.sv:20:5
						VX_reset_relay #(
							.N(1),
							.MAX_FANOUT(0)
						) __icache_reset(
							.clk(clk),
							.reset(reset),
							.reset_o(icache_reset)
						);
						// Trace: src/VX_socket.sv:25:5
						// expanded module instance: icache
						localparam _bbase_9B047_core_bus_if = 0;
						localparam _bbase_9B047_mem_bus_if = 0;
						localparam _param_9B047_INSTANCE_ID = "";
						localparam _param_9B047_NUM_UNITS = 1;
						localparam _param_9B047_NUM_INPUTS = 1;
						localparam _param_9B047_TAG_SEL_IDX = 0;
						localparam _param_9B047_CACHE_SIZE = 16384;
						localparam _param_9B047_LINE_SIZE = VX_gpu_pkg_ICACHE_LINE_SIZE;
						localparam _param_9B047_NUM_BANKS = 1;
						localparam _param_9B047_NUM_WAYS = 4;
						localparam _param_9B047_WORD_SIZE = VX_gpu_pkg_ICACHE_WORD_SIZE;
						localparam _param_9B047_NUM_REQS = 1;
						localparam _param_9B047_MEM_PORTS = 1;
						localparam _param_9B047_CRSQ_SIZE = 2;
						localparam _param_9B047_MSHR_SIZE = 16;
						localparam _param_9B047_MRSQ_SIZE = 0;
						localparam _param_9B047_MREQ_SIZE = 4;
						localparam _param_9B047_TAG_WIDTH = VX_gpu_pkg_ICACHE_TAG_WIDTH;
						localparam _param_9B047_WRITE_ENABLE = 0;
						localparam _param_9B047_REPL_POLICY = 1;
						localparam _param_9B047_NC_ENABLE = 0;
						localparam _param_9B047_CORE_OUT_BUF = 3;
						localparam _param_9B047_MEM_OUT_BUF = 2;
						if (1) begin : icache
							// removed import VX_gpu_pkg::*;
							// Trace: src/VX_cache_cluster.sv:2:15
							localparam INSTANCE_ID = _param_9B047_INSTANCE_ID;
							// Trace: src/VX_cache_cluster.sv:3:15
							localparam NUM_UNITS = _param_9B047_NUM_UNITS;
							// Trace: src/VX_cache_cluster.sv:4:15
							localparam NUM_INPUTS = _param_9B047_NUM_INPUTS;
							// Trace: src/VX_cache_cluster.sv:5:15
							localparam TAG_SEL_IDX = _param_9B047_TAG_SEL_IDX;
							// Trace: src/VX_cache_cluster.sv:6:15
							localparam NUM_REQS = _param_9B047_NUM_REQS;
							// Trace: src/VX_cache_cluster.sv:7:15
							localparam MEM_PORTS = _param_9B047_MEM_PORTS;
							// Trace: src/VX_cache_cluster.sv:8:15
							localparam CACHE_SIZE = _param_9B047_CACHE_SIZE;
							// Trace: src/VX_cache_cluster.sv:9:15
							localparam LINE_SIZE = _param_9B047_LINE_SIZE;
							// Trace: src/VX_cache_cluster.sv:10:15
							localparam NUM_BANKS = _param_9B047_NUM_BANKS;
							// Trace: src/VX_cache_cluster.sv:11:15
							localparam NUM_WAYS = _param_9B047_NUM_WAYS;
							// Trace: src/VX_cache_cluster.sv:12:15
							localparam WORD_SIZE = _param_9B047_WORD_SIZE;
							// Trace: src/VX_cache_cluster.sv:13:15
							localparam CRSQ_SIZE = _param_9B047_CRSQ_SIZE;
							// Trace: src/VX_cache_cluster.sv:14:15
							localparam MSHR_SIZE = _param_9B047_MSHR_SIZE;
							// Trace: src/VX_cache_cluster.sv:15:15
							localparam MRSQ_SIZE = _param_9B047_MRSQ_SIZE;
							// Trace: src/VX_cache_cluster.sv:16:15
							localparam MREQ_SIZE = _param_9B047_MREQ_SIZE;
							// Trace: src/VX_cache_cluster.sv:17:15
							localparam WRITE_ENABLE = _param_9B047_WRITE_ENABLE;
							// Trace: src/VX_cache_cluster.sv:18:15
							localparam WRITEBACK = 0;
							// Trace: src/VX_cache_cluster.sv:19:15
							localparam DIRTY_BYTES = 0;
							// Trace: src/VX_cache_cluster.sv:20:15
							localparam REPL_POLICY = _param_9B047_REPL_POLICY;
							// Trace: src/VX_cache_cluster.sv:21:15
							localparam VX_gpu_pkg_UUID_WIDTH = 1;
							localparam TAG_WIDTH = _param_9B047_TAG_WIDTH;
							// Trace: src/VX_cache_cluster.sv:22:15
							localparam NC_ENABLE = _param_9B047_NC_ENABLE;
							// Trace: src/VX_cache_cluster.sv:23:15
							localparam CORE_OUT_BUF = _param_9B047_CORE_OUT_BUF;
							// Trace: src/VX_cache_cluster.sv:24:15
							localparam MEM_OUT_BUF = _param_9B047_MEM_OUT_BUF;
							// Trace: src/VX_cache_cluster.sv:26:5
							wire clk;
							// Trace: src/VX_cache_cluster.sv:27:5
							wire reset;
							// Trace: src/VX_cache_cluster.sv:28:5
							localparam _mbase_core_bus_if = 0;
							// Trace: src/VX_cache_cluster.sv:29:5
							localparam _mbase_mem_bus_if = 0;
							// Trace: src/VX_cache_cluster.sv:31:5
							localparam NUM_CACHES = NUM_UNITS;
							// Trace: src/VX_cache_cluster.sv:32:5
							localparam PASSTHRU = 1'd0;
							// Trace: src/VX_cache_cluster.sv:33:5
							localparam ARB_TAG_WIDTH = 3;
							// Trace: src/VX_cache_cluster.sv:34:5
							localparam CACHE_MEM_TAG_WIDTH = 5;
							// Trace: src/VX_cache_cluster.sv:36:5
							localparam BYPASS_TAG_WIDTH = 7;
							// Trace: src/VX_cache_cluster.sv:38:5
							localparam NC_TAG_WIDTH = 8;
							// Trace: src/VX_cache_cluster.sv:39:5
							localparam MEM_TAG_WIDTH = (PASSTHRU ? BYPASS_TAG_WIDTH : (NC_ENABLE ? NC_TAG_WIDTH : CACHE_MEM_TAG_WIDTH));
							// Trace: src/VX_cache_cluster.sv:40:5
							// expanded interface instance: cache_mem_bus_if
							localparam _param_A4879_DATA_SIZE = LINE_SIZE;
							localparam _param_A4879_TAG_WIDTH = MEM_TAG_WIDTH;
							genvar _arr_A4879;
							for (_arr_A4879 = 0; _arr_A4879 <= 0; _arr_A4879 = _arr_A4879 + 1) begin : cache_mem_bus_if
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_A4879_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
								localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
								localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_A4879_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:8:5
								localparam VX_gpu_pkg_UUID_WIDTH = 1;
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:12:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:20:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:24:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire [610:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire [516:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:30:5
								// Trace: src/VX_mem_bus_if.sv:38:5
							end
							// Trace: src/VX_cache_cluster.sv:44:5
							// expanded interface instance: arb_core_bus_if
							localparam _param_F9BC9_DATA_SIZE = WORD_SIZE;
							localparam _param_F9BC9_TAG_WIDTH = ARB_TAG_WIDTH;
							genvar _arr_F9BC9;
							for (_arr_F9BC9 = 0; _arr_F9BC9 <= 0; _arr_F9BC9 = _arr_F9BC9 + 1) begin : arb_core_bus_if
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_F9BC9_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
								localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
								localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_F9BC9_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 30;
								// Trace: src/VX_mem_bus_if.sv:8:5
								localparam VX_gpu_pkg_UUID_WIDTH = 1;
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:12:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:20:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:24:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire [72:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire [34:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:30:5
								// Trace: src/VX_mem_bus_if.sv:38:5
							end
							// Trace: src/VX_cache_cluster.sv:48:5
							genvar _gv_i_191;
							for (_gv_i_191 = 0; _gv_i_191 < NUM_REQS; _gv_i_191 = _gv_i_191 + 1) begin : g_core_arb
								localparam i = _gv_i_191;
								// Trace: src/VX_cache_cluster.sv:49:9
								// expanded interface instance: core_bus_tmp_if
								localparam _param_A62F7_DATA_SIZE = WORD_SIZE;
								localparam _param_A62F7_TAG_WIDTH = TAG_WIDTH;
								genvar _arr_A62F7;
								for (_arr_A62F7 = 0; _arr_A62F7 <= 0; _arr_A62F7 = _arr_A62F7 + 1) begin : core_bus_tmp_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_A62F7_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_A62F7_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 30;
									// Trace: src/VX_mem_bus_if.sv:8:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:12:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:20:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:24:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire [72:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire [34:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:30:5
									// Trace: src/VX_mem_bus_if.sv:38:5
								end
								// Trace: src/VX_cache_cluster.sv:53:9
								// expanded interface instance: arb_core_bus_tmp_if
								localparam _param_E788B_DATA_SIZE = WORD_SIZE;
								localparam _param_E788B_TAG_WIDTH = ARB_TAG_WIDTH;
								genvar _arr_E788B;
								for (_arr_E788B = 0; _arr_E788B <= 0; _arr_E788B = _arr_E788B + 1) begin : arb_core_bus_tmp_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_E788B_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_E788B_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 30;
									// Trace: src/VX_mem_bus_if.sv:8:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:12:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:20:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:24:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire [72:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire [34:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:30:5
									// Trace: src/VX_mem_bus_if.sv:38:5
								end
								genvar _gv_j_19;
								for (_gv_j_19 = 0; _gv_j_19 < NUM_INPUTS; _gv_j_19 = _gv_j_19 + 1) begin : g_core_bus_tmp_if
									localparam j = _gv_j_19;
									// Trace: src/VX_cache_cluster.sv:58:5
									assign core_bus_tmp_if[j].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].req_valid;
									// Trace: src/VX_cache_cluster.sv:59:5
									assign core_bus_tmp_if[j].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].req_data;
									// Trace: src/VX_cache_cluster.sv:60:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].req_ready = core_bus_tmp_if[j].req_ready;
									// Trace: src/VX_cache_cluster.sv:61:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].rsp_valid = core_bus_tmp_if[j].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:62:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].rsp_data = core_bus_tmp_if[j].rsp_data;
									// Trace: src/VX_cache_cluster.sv:63:5
									assign core_bus_tmp_if[j].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].rsp_ready;
								end
								// Trace: src/VX_cache_cluster.sv:65:9
								// expanded module instance: core_arb
								localparam _bbase_856A9_bus_in_if = 0;
								localparam _bbase_856A9_bus_out_if = 0;
								localparam _param_856A9_NUM_INPUTS = NUM_INPUTS;
								localparam _param_856A9_NUM_OUTPUTS = NUM_CACHES;
								localparam _param_856A9_DATA_SIZE = WORD_SIZE;
								localparam _param_856A9_TAG_WIDTH = TAG_WIDTH;
								localparam _param_856A9_TAG_SEL_IDX = TAG_SEL_IDX;
								localparam _param_856A9_ARBITER = "R";
								localparam _param_856A9_REQ_OUT_BUF = 0;
								localparam _param_856A9_RSP_OUT_BUF = 0;
								if (1) begin : core_arb
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_arb.sv:2:15
									localparam NUM_INPUTS = _param_856A9_NUM_INPUTS;
									// Trace: src/VX_mem_arb.sv:3:15
									localparam NUM_OUTPUTS = _param_856A9_NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:4:15
									localparam DATA_SIZE = _param_856A9_DATA_SIZE;
									// Trace: src/VX_mem_arb.sv:5:15
									localparam TAG_WIDTH = _param_856A9_TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:6:15
									localparam TAG_SEL_IDX = _param_856A9_TAG_SEL_IDX;
									// Trace: src/VX_mem_arb.sv:7:15
									localparam REQ_OUT_BUF = _param_856A9_REQ_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:8:15
									localparam RSP_OUT_BUF = _param_856A9_RSP_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:9:15
									localparam ARBITER = _param_856A9_ARBITER;
									// Trace: src/VX_mem_arb.sv:10:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_arb.sv:11:15
									localparam ADDR_WIDTH = 30;
									// Trace: src/VX_mem_arb.sv:12:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_arb.sv:14:5
									wire clk;
									// Trace: src/VX_mem_arb.sv:15:5
									wire reset;
									// Trace: src/VX_mem_arb.sv:16:5
									localparam _mbase_bus_in_if = 0;
									// Trace: src/VX_mem_arb.sv:17:5
									localparam _mbase_bus_out_if = 0;
									// Trace: src/VX_mem_arb.sv:19:5
									localparam DATA_WIDTH = 32;
									// Trace: src/VX_mem_arb.sv:20:5
									localparam LOG_NUM_REQS = 0;
									// Trace: src/VX_mem_arb.sv:21:5
									localparam REQ_DATAW = 73;
									// Trace: src/VX_mem_arb.sv:22:5
									localparam RSP_DATAW = 35;
									// Trace: src/VX_mem_arb.sv:23:5
									localparam SEL_COUNT = NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:24:5
									wire [0:0] req_valid_in;
									// Trace: src/VX_mem_arb.sv:25:5
									wire [72:0] req_data_in;
									// Trace: src/VX_mem_arb.sv:26:5
									wire [0:0] req_ready_in;
									// Trace: src/VX_mem_arb.sv:27:5
									wire [0:0] req_valid_out;
									// Trace: src/VX_mem_arb.sv:28:5
									wire [72:0] req_data_out;
									// Trace: src/VX_mem_arb.sv:29:5
									wire [0:0] req_sel_out;
									// Trace: src/VX_mem_arb.sv:30:5
									wire [0:0] req_ready_out;
									// Trace: src/VX_mem_arb.sv:31:5
									genvar _gv_i_183;
									for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
										localparam i = _gv_i_183;
										// Trace: src/VX_mem_arb.sv:32:9
										assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].core_bus_tmp_if[i + _mbase_bus_in_if].req_valid;
										// Trace: src/VX_mem_arb.sv:33:9
										assign req_data_in[i * 73+:73] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].core_bus_tmp_if[i + _mbase_bus_in_if].req_data;
										// Trace: src/VX_mem_arb.sv:34:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].core_bus_tmp_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:36:5
									VX_stream_arb #(
										.NUM_INPUTS(NUM_INPUTS),
										.NUM_OUTPUTS(NUM_OUTPUTS),
										.DATAW(REQ_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(REQ_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(req_valid_in),
										.ready_in(req_ready_in),
										.data_in(req_data_in),
										.data_out(req_data_out),
										.sel_out(req_sel_out),
										.valid_out(req_valid_out),
										.ready_out(req_ready_out)
									);
									// Trace: src/VX_mem_arb.sv:53:5
									genvar _gv_i_184;
									for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
										localparam i = _gv_i_184;
										// Trace: src/VX_mem_arb.sv:54:9
										wire [2:0] req_tag_out;
										// Trace: src/VX_mem_arb.sv:55:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
										// Trace: src/VX_mem_arb.sv:56:9
										assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[72], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[71-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[41-:32], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[9-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[5-:3], req_tag_out} = req_data_out[i * 73+:73];
										// Trace: src/VX_mem_arb.sv:64:9
										assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
										if (1) begin : g_req_tag_out
											// Trace: src/VX_mem_arb.sv:76:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[2-:3] = req_tag_out;
										end
									end
									// Trace: src/VX_mem_arb.sv:79:5
									wire [0:0] rsp_valid_out;
									// Trace: src/VX_mem_arb.sv:80:5
									wire [34:0] rsp_data_out;
									// Trace: src/VX_mem_arb.sv:81:5
									wire [0:0] rsp_ready_out;
									// Trace: src/VX_mem_arb.sv:82:5
									wire [0:0] rsp_valid_in;
									// Trace: src/VX_mem_arb.sv:83:5
									wire [34:0] rsp_data_in;
									// Trace: src/VX_mem_arb.sv:84:5
									wire [0:0] rsp_ready_in;
									// Trace: src/VX_mem_arb.sv:85:5
									if (1) begin : g_rsp_arb
										genvar _gv_i_186;
										for (_gv_i_186 = 0; _gv_i_186 < NUM_OUTPUTS; _gv_i_186 = _gv_i_186 + 1) begin : g_rsp_data_in
											localparam i = _gv_i_186;
											// Trace: src/VX_mem_arb.sv:120:13
											assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
											// Trace: src/VX_mem_arb.sv:121:13
											assign rsp_data_in[i * 35+:35] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
											// Trace: src/VX_mem_arb.sv:122:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
										end
										// Trace: src/VX_mem_arb.sv:124:9
										VX_stream_arb #(
											.NUM_INPUTS(NUM_OUTPUTS),
											.NUM_OUTPUTS(NUM_INPUTS),
											.DATAW(RSP_DATAW),
											.ARBITER(ARBITER),
											.OUT_BUF(RSP_OUT_BUF)
										) req_arb(
											.clk(clk),
											.reset(reset),
											.valid_in(rsp_valid_in),
											.ready_in(rsp_ready_in),
											.data_in(rsp_data_in),
											.data_out(rsp_data_out),
											.valid_out(rsp_valid_out),
											.ready_out(rsp_ready_out),
											.sel_out()
										);
									end
									// Trace: src/VX_mem_arb.sv:142:5
									genvar _gv_i_187;
									for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
										localparam i = _gv_i_187;
										// Trace: src/VX_mem_arb.sv:143:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].core_bus_tmp_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
										// Trace: src/VX_mem_arb.sv:144:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].core_bus_tmp_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 35+:35];
										// Trace: src/VX_mem_arb.sv:145:9
										assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_core_arb[_gv_i_191].core_bus_tmp_if[i + _mbase_bus_in_if].rsp_ready;
									end
								end
								assign core_arb.clk = clk;
								assign core_arb.reset = reset;
								genvar _gv_k_1;
								for (_gv_k_1 = 0; _gv_k_1 < NUM_CACHES; _gv_k_1 = _gv_k_1 + 1) begin : g_arb_core_bus_if
									localparam k = _gv_k_1;
									// Trace: src/VX_cache_cluster.sv:81:5
									assign arb_core_bus_if[(k * NUM_REQS) + i].req_valid = arb_core_bus_tmp_if[k].req_valid;
									// Trace: src/VX_cache_cluster.sv:82:5
									assign arb_core_bus_if[(k * NUM_REQS) + i].req_data = arb_core_bus_tmp_if[k].req_data;
									// Trace: src/VX_cache_cluster.sv:83:5
									assign arb_core_bus_tmp_if[k].req_ready = arb_core_bus_if[(k * NUM_REQS) + i].req_ready;
									// Trace: src/VX_cache_cluster.sv:84:5
									assign arb_core_bus_tmp_if[k].rsp_valid = arb_core_bus_if[(k * NUM_REQS) + i].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:85:5
									assign arb_core_bus_tmp_if[k].rsp_data = arb_core_bus_if[(k * NUM_REQS) + i].rsp_data;
									// Trace: src/VX_cache_cluster.sv:86:5
									assign arb_core_bus_if[(k * NUM_REQS) + i].rsp_ready = arb_core_bus_tmp_if[k].rsp_ready;
								end
							end
							// Trace: src/VX_cache_cluster.sv:89:6
							genvar _gv_i_192;
							for (_gv_i_192 = 0; _gv_i_192 < NUM_CACHES; _gv_i_192 = _gv_i_192 + 1) begin : g_cache_wrap
								localparam i = _gv_i_192;
								// Trace: src/VX_cache_cluster.sv:90:9
								// expanded module instance: cache_wrap
								localparam _bbase_665FE_core_bus_if = i * NUM_REQS;
								localparam _bbase_665FE_mem_bus_if = i * MEM_PORTS;
								localparam _param_665FE_INSTANCE_ID = "";
								localparam _param_665FE_CACHE_SIZE = CACHE_SIZE;
								localparam _param_665FE_LINE_SIZE = LINE_SIZE;
								localparam _param_665FE_NUM_BANKS = NUM_BANKS;
								localparam _param_665FE_NUM_WAYS = NUM_WAYS;
								localparam _param_665FE_WORD_SIZE = WORD_SIZE;
								localparam _param_665FE_NUM_REQS = NUM_REQS;
								localparam _param_665FE_MEM_PORTS = MEM_PORTS;
								localparam _param_665FE_WRITE_ENABLE = WRITE_ENABLE;
								localparam _param_665FE_WRITEBACK = WRITEBACK;
								localparam _param_665FE_DIRTY_BYTES = DIRTY_BYTES;
								localparam _param_665FE_REPL_POLICY = REPL_POLICY;
								localparam _param_665FE_CRSQ_SIZE = CRSQ_SIZE;
								localparam _param_665FE_MSHR_SIZE = MSHR_SIZE;
								localparam _param_665FE_MRSQ_SIZE = MRSQ_SIZE;
								localparam _param_665FE_MREQ_SIZE = MREQ_SIZE;
								localparam _param_665FE_TAG_WIDTH = ARB_TAG_WIDTH;
								localparam _param_665FE_TAG_SEL_IDX = TAG_SEL_IDX;
								localparam _param_665FE_CORE_OUT_BUF = CORE_OUT_BUF;
								localparam _param_665FE_MEM_OUT_BUF = MEM_OUT_BUF;
								localparam _param_665FE_NC_ENABLE = NC_ENABLE;
								localparam _param_665FE_PASSTHRU = PASSTHRU;
								if (1) begin : cache_wrap
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_cache_wrap.sv:2:15
									localparam INSTANCE_ID = _param_665FE_INSTANCE_ID;
									// Trace: src/VX_cache_wrap.sv:3:15
									localparam TAG_SEL_IDX = _param_665FE_TAG_SEL_IDX;
									// Trace: src/VX_cache_wrap.sv:4:15
									localparam NUM_REQS = _param_665FE_NUM_REQS;
									// Trace: src/VX_cache_wrap.sv:5:15
									localparam MEM_PORTS = _param_665FE_MEM_PORTS;
									// Trace: src/VX_cache_wrap.sv:6:15
									localparam CACHE_SIZE = _param_665FE_CACHE_SIZE;
									// Trace: src/VX_cache_wrap.sv:7:15
									localparam LINE_SIZE = _param_665FE_LINE_SIZE;
									// Trace: src/VX_cache_wrap.sv:8:15
									localparam NUM_BANKS = _param_665FE_NUM_BANKS;
									// Trace: src/VX_cache_wrap.sv:9:15
									localparam NUM_WAYS = _param_665FE_NUM_WAYS;
									// Trace: src/VX_cache_wrap.sv:10:15
									localparam WORD_SIZE = _param_665FE_WORD_SIZE;
									// Trace: src/VX_cache_wrap.sv:11:15
									localparam CRSQ_SIZE = _param_665FE_CRSQ_SIZE;
									// Trace: src/VX_cache_wrap.sv:12:15
									localparam MSHR_SIZE = _param_665FE_MSHR_SIZE;
									// Trace: src/VX_cache_wrap.sv:13:15
									localparam MRSQ_SIZE = _param_665FE_MRSQ_SIZE;
									// Trace: src/VX_cache_wrap.sv:14:15
									localparam MREQ_SIZE = _param_665FE_MREQ_SIZE;
									// Trace: src/VX_cache_wrap.sv:15:15
									localparam WRITE_ENABLE = _param_665FE_WRITE_ENABLE;
									// Trace: src/VX_cache_wrap.sv:16:15
									localparam WRITEBACK = _param_665FE_WRITEBACK;
									// Trace: src/VX_cache_wrap.sv:17:15
									localparam DIRTY_BYTES = _param_665FE_DIRTY_BYTES;
									// Trace: src/VX_cache_wrap.sv:18:15
									localparam REPL_POLICY = _param_665FE_REPL_POLICY;
									// Trace: src/VX_cache_wrap.sv:19:15
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									localparam TAG_WIDTH = _param_665FE_TAG_WIDTH;
									// Trace: src/VX_cache_wrap.sv:20:15
									localparam NC_ENABLE = _param_665FE_NC_ENABLE;
									// Trace: src/VX_cache_wrap.sv:21:15
									localparam PASSTHRU = _param_665FE_PASSTHRU;
									// Trace: src/VX_cache_wrap.sv:22:15
									localparam CORE_OUT_BUF = _param_665FE_CORE_OUT_BUF;
									// Trace: src/VX_cache_wrap.sv:23:15
									localparam MEM_OUT_BUF = _param_665FE_MEM_OUT_BUF;
									// Trace: src/VX_cache_wrap.sv:25:5
									wire clk;
									// Trace: src/VX_cache_wrap.sv:26:5
									wire reset;
									// Trace: src/VX_cache_wrap.sv:27:5
									localparam _mbase_core_bus_if = _bbase_665FE_core_bus_if;
									// Trace: src/VX_cache_wrap.sv:28:5
									localparam _mbase_mem_bus_if = _bbase_665FE_mem_bus_if;
									// Trace: src/VX_cache_wrap.sv:30:5
									localparam CACHE_MEM_TAG_WIDTH = 5;
									// Trace: src/VX_cache_wrap.sv:32:5
									localparam BYPASS_TAG_WIDTH = 7;
									// Trace: src/VX_cache_wrap.sv:34:5
									localparam NC_TAG_WIDTH = 8;
									// Trace: src/VX_cache_wrap.sv:35:5
									localparam MEM_TAG_WIDTH = (PASSTHRU ? BYPASS_TAG_WIDTH : (NC_ENABLE ? NC_TAG_WIDTH : CACHE_MEM_TAG_WIDTH));
									// Trace: src/VX_cache_wrap.sv:36:5
									localparam BYPASS_ENABLE = 1'd0;
									// Trace: src/VX_cache_wrap.sv:37:5
									// expanded interface instance: core_bus_cache_if
									localparam _param_24C1C_DATA_SIZE = WORD_SIZE;
									localparam _param_24C1C_TAG_WIDTH = TAG_WIDTH;
									genvar _arr_24C1C;
									for (_arr_24C1C = 0; _arr_24C1C <= 0; _arr_24C1C = _arr_24C1C + 1) begin : core_bus_cache_if
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_24C1C_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_24C1C_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 30;
										// Trace: src/VX_mem_bus_if.sv:8:5
										localparam VX_gpu_pkg_UUID_WIDTH = 1;
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:12:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:20:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:24:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire [72:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire [34:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:30:5
										// Trace: src/VX_mem_bus_if.sv:38:5
									end
									// Trace: src/VX_cache_wrap.sv:41:5
									// expanded interface instance: mem_bus_cache_if
									localparam _param_D895D_DATA_SIZE = LINE_SIZE;
									localparam _param_D895D_TAG_WIDTH = CACHE_MEM_TAG_WIDTH;
									genvar _arr_D895D;
									for (_arr_D895D = 0; _arr_D895D <= 0; _arr_D895D = _arr_D895D + 1) begin : mem_bus_cache_if
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_D895D_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_D895D_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 26;
										// Trace: src/VX_mem_bus_if.sv:8:5
										localparam VX_gpu_pkg_UUID_WIDTH = 1;
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:12:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:20:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:24:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire [610:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire [516:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:30:5
										// Trace: src/VX_mem_bus_if.sv:38:5
									end
									// Trace: src/VX_cache_wrap.sv:45:5
									// expanded interface instance: mem_bus_tmp_if
									localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
									localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH;
									genvar _arr_4FE36;
									for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 26;
										// Trace: src/VX_mem_bus_if.sv:8:5
										localparam VX_gpu_pkg_UUID_WIDTH = 1;
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:12:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:20:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:24:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire [610:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire [516:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:30:5
										// Trace: src/VX_mem_bus_if.sv:38:5
									end
									// Trace: src/VX_cache_wrap.sv:49:5
									if (BYPASS_ENABLE) begin : g_bypass
										// Trace: src/VX_cache_wrap.sv:50:9
										// expanded module instance: cache_bypass
										localparam _bbase_714AA_core_bus_in_if = i * NUM_REQS;
										localparam _bbase_714AA_core_bus_out_if = 0;
										localparam _bbase_714AA_mem_bus_in_if = 0;
										localparam _bbase_714AA_mem_bus_out_if = 0;
										localparam _param_714AA_NUM_REQS = NUM_REQS;
										localparam _param_714AA_MEM_PORTS = MEM_PORTS;
										localparam _param_714AA_TAG_SEL_IDX = TAG_SEL_IDX;
										localparam _param_714AA_CACHE_ENABLE = !PASSTHRU;
										localparam _param_714AA_WORD_SIZE = WORD_SIZE;
										localparam _param_714AA_LINE_SIZE = LINE_SIZE;
										localparam _param_714AA_CORE_ADDR_WIDTH = 30;
										localparam _param_714AA_CORE_TAG_WIDTH = TAG_WIDTH;
										localparam _param_714AA_MEM_ADDR_WIDTH = 26;
										localparam _param_714AA_MEM_TAG_IN_WIDTH = CACHE_MEM_TAG_WIDTH;
										localparam _param_714AA_CORE_OUT_BUF = CORE_OUT_BUF;
										localparam _param_714AA_MEM_OUT_BUF = MEM_OUT_BUF;
										if (1) begin : cache_bypass
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_cache_bypass.sv:2:15
											localparam NUM_REQS = _param_714AA_NUM_REQS;
											// Trace: src/VX_cache_bypass.sv:3:15
											localparam MEM_PORTS = _param_714AA_MEM_PORTS;
											// Trace: src/VX_cache_bypass.sv:4:15
											localparam TAG_SEL_IDX = _param_714AA_TAG_SEL_IDX;
											// Trace: src/VX_cache_bypass.sv:5:15
											localparam CACHE_ENABLE = _param_714AA_CACHE_ENABLE;
											// Trace: src/VX_cache_bypass.sv:6:15
											localparam WORD_SIZE = _param_714AA_WORD_SIZE;
											// Trace: src/VX_cache_bypass.sv:7:15
											localparam LINE_SIZE = _param_714AA_LINE_SIZE;
											// Trace: src/VX_cache_bypass.sv:8:15
											localparam CORE_ADDR_WIDTH = _param_714AA_CORE_ADDR_WIDTH;
											// Trace: src/VX_cache_bypass.sv:9:15
											localparam CORE_TAG_WIDTH = _param_714AA_CORE_TAG_WIDTH;
											// Trace: src/VX_cache_bypass.sv:10:15
											localparam MEM_ADDR_WIDTH = _param_714AA_MEM_ADDR_WIDTH;
											// Trace: src/VX_cache_bypass.sv:11:15
											localparam MEM_TAG_IN_WIDTH = _param_714AA_MEM_TAG_IN_WIDTH;
											// Trace: src/VX_cache_bypass.sv:12:15
											localparam CORE_OUT_BUF = _param_714AA_CORE_OUT_BUF;
											// Trace: src/VX_cache_bypass.sv:13:15
											localparam MEM_OUT_BUF = _param_714AA_MEM_OUT_BUF;
											// Trace: src/VX_cache_bypass.sv:15:5
											wire clk;
											// Trace: src/VX_cache_bypass.sv:16:5
											wire reset;
											// Trace: src/VX_cache_bypass.sv:17:5
											localparam _mbase_core_bus_in_if = _bbase_714AA_core_bus_in_if;
											// Trace: src/VX_cache_bypass.sv:18:5
											localparam _mbase_core_bus_out_if = 0;
											// Trace: src/VX_cache_bypass.sv:19:5
											localparam _mbase_mem_bus_in_if = 0;
											// Trace: src/VX_cache_bypass.sv:20:5
											localparam _mbase_mem_bus_out_if = 0;
											// Trace: src/VX_cache_bypass.sv:22:5
											localparam DIRECT_PASSTHRU = (!CACHE_ENABLE && 1'd0) && 1'd1;
											// Trace: src/VX_cache_bypass.sv:23:5
											localparam CORE_DATA_WIDTH = 32;
											// Trace: src/VX_cache_bypass.sv:24:5
											localparam WORDS_PER_LINE = 16;
											// Trace: src/VX_cache_bypass.sv:25:5
											localparam WSEL_BITS = 4;
											// Trace: src/VX_cache_bypass.sv:26:5
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam CORE_TAG_ID_WIDTH = 2;
											// Trace: src/VX_cache_bypass.sv:27:5
											localparam MEM_TAG_ID_WIDTH = 2;
											// Trace: src/VX_cache_bypass.sv:28:5
											localparam MEM_TAG_NC1_WIDTH = 3;
											// Trace: src/VX_cache_bypass.sv:29:5
											localparam MEM_TAG_NC2_WIDTH = 7;
											// Trace: src/VX_cache_bypass.sv:30:5
											localparam MEM_TAG_OUT_WIDTH = (CACHE_ENABLE ? MEM_TAG_NC2_WIDTH : MEM_TAG_NC2_WIDTH);
											// Trace: src/VX_cache_bypass.sv:31:5
											// expanded interface instance: core_bus_nc_switch_if
											localparam _param_95306_DATA_SIZE = WORD_SIZE;
											localparam _param_95306_TAG_WIDTH = CORE_TAG_WIDTH;
											genvar _arr_95306;
											for (_arr_95306 = 0; _arr_95306 <= (((CACHE_ENABLE ? 2 : 1) * NUM_REQS) - 1); _arr_95306 = _arr_95306 + 1) begin : core_bus_nc_switch_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_95306_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_95306_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 30;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [72:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [34:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache_bypass.sv:35:5
											wire [0:0] core_req_nc_sel;
											// Trace: src/VX_cache_bypass.sv:36:5
											genvar _gv_i_56;
											localparam VX_gpu_pkg_MEM_REQ_FLAG_IO = 1;
											for (_gv_i_56 = 0; _gv_i_56 < NUM_REQS; _gv_i_56 = _gv_i_56 + 1) begin : g_core_req_is_nc
												localparam i = _gv_i_56;
												if (CACHE_ENABLE) begin : g_cache
													// Trace: src/VX_cache_bypass.sv:38:13
													assign core_req_nc_sel[i] = ~Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_in_if].req_data[4];
												end
												else begin : g_no_cache
													// Trace: src/VX_cache_bypass.sv:40:13
													assign core_req_nc_sel[i] = 1'b0;
												end
											end
											// Trace: src/VX_cache_bypass.sv:43:5
											// expanded module instance: core_bus_nc_switch
											localparam _bbase_69FDB_bus_in_if = i * NUM_REQS;
											localparam _bbase_69FDB_bus_out_if = 0;
											localparam _param_69FDB_NUM_INPUTS = NUM_REQS;
											localparam _param_69FDB_NUM_OUTPUTS = (CACHE_ENABLE ? 2 : 1) * NUM_REQS;
											localparam _param_69FDB_DATA_SIZE = WORD_SIZE;
											localparam _param_69FDB_TAG_WIDTH = CORE_TAG_WIDTH;
											localparam _param_69FDB_ARBITER = "R";
											localparam _param_69FDB_REQ_OUT_BUF = 0;
											localparam _param_69FDB_RSP_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
											if (1) begin : core_bus_nc_switch
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_switch.sv:2:15
												localparam NUM_INPUTS = _param_69FDB_NUM_INPUTS;
												// Trace: src/VX_mem_switch.sv:3:15
												localparam NUM_OUTPUTS = _param_69FDB_NUM_OUTPUTS;
												// Trace: src/VX_mem_switch.sv:4:15
												localparam DATA_SIZE = _param_69FDB_DATA_SIZE;
												// Trace: src/VX_mem_switch.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_switch.sv:6:15
												localparam ADDR_WIDTH = 30;
												// Trace: src/VX_mem_switch.sv:7:15
												localparam TAG_WIDTH = _param_69FDB_TAG_WIDTH;
												// Trace: src/VX_mem_switch.sv:8:15
												localparam REQ_OUT_BUF = _param_69FDB_REQ_OUT_BUF;
												// Trace: src/VX_mem_switch.sv:9:15
												localparam RSP_OUT_BUF = _param_69FDB_RSP_OUT_BUF;
												// Trace: src/VX_mem_switch.sv:10:15
												localparam ARBITER = _param_69FDB_ARBITER;
												// Trace: src/VX_mem_switch.sv:11:15
												localparam NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? ((NUM_INPUTS + NUM_OUTPUTS) - 1) / NUM_OUTPUTS : ((NUM_OUTPUTS + NUM_INPUTS) - 1) / NUM_INPUTS);
												// Trace: src/VX_mem_switch.sv:12:15
												localparam SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
												// Trace: src/VX_mem_switch.sv:13:15
												localparam LOG_NUM_REQS = $clog2(NUM_REQS);
												// Trace: src/VX_mem_switch.sv:15:5
												wire clk;
												// Trace: src/VX_mem_switch.sv:16:5
												wire reset;
												// Trace: src/VX_mem_switch.sv:17:5
												wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] bus_sel;
												// Trace: src/VX_mem_switch.sv:18:5
												localparam _mbase_bus_in_if = _bbase_69FDB_bus_in_if;
												// Trace: src/VX_mem_switch.sv:19:5
												localparam _mbase_bus_out_if = 0;
												// Trace: src/VX_mem_switch.sv:21:5
												localparam DATA_WIDTH = 32;
												// Trace: src/VX_mem_switch.sv:22:5
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam REQ_DATAW = 73;
												// Trace: src/VX_mem_switch.sv:23:5
												localparam RSP_DATAW = 35;
												// Trace: src/VX_mem_switch.sv:24:5
												wire [0:0] req_valid_in;
												// Trace: src/VX_mem_switch.sv:25:5
												wire [72:0] req_data_in;
												// Trace: src/VX_mem_switch.sv:26:5
												wire [0:0] req_ready_in;
												// Trace: src/VX_mem_switch.sv:27:5
												wire [NUM_OUTPUTS - 1:0] req_valid_out;
												// Trace: src/VX_mem_switch.sv:28:5
												wire [(NUM_OUTPUTS * 73) - 1:0] req_data_out;
												// Trace: src/VX_mem_switch.sv:29:5
												wire [NUM_OUTPUTS - 1:0] req_ready_out;
												// Trace: src/VX_mem_switch.sv:30:5
												genvar _gv_i_109;
												for (_gv_i_109 = 0; _gv_i_109 < NUM_INPUTS; _gv_i_109 = _gv_i_109 + 1) begin : g_req_data_in
													localparam i = _gv_i_109;
													// Trace: src/VX_mem_switch.sv:31:9
													assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_bus_in_if].req_valid;
													// Trace: src/VX_mem_switch.sv:32:9
													assign req_data_in[i * 73+:73] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_bus_in_if].req_data;
													// Trace: src/VX_mem_switch.sv:33:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
												end
												// Trace: src/VX_mem_switch.sv:35:5
												VX_stream_switch #(
													.NUM_INPUTS(NUM_INPUTS),
													.NUM_OUTPUTS(NUM_OUTPUTS),
													.DATAW(REQ_DATAW),
													.OUT_BUF(REQ_OUT_BUF)
												) req_switch(
													.clk(clk),
													.reset(reset),
													.sel_in(bus_sel),
													.valid_in(req_valid_in),
													.data_in(req_data_in),
													.ready_in(req_ready_in),
													.valid_out(req_valid_out),
													.data_out(req_data_out),
													.ready_out(req_ready_out)
												);
												// Trace: src/VX_mem_switch.sv:51:5
												genvar _gv_i_110;
												for (_gv_i_110 = 0; _gv_i_110 < NUM_OUTPUTS; _gv_i_110 = _gv_i_110 + 1) begin : g_req_data_out
													localparam i = _gv_i_110;
													// Trace: src/VX_mem_switch.sv:52:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
													// Trace: src/VX_mem_switch.sv:53:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_data = req_data_out[i * 73+:73];
													// Trace: src/VX_mem_switch.sv:54:9
													assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_ready;
												end
												// Trace: src/VX_mem_switch.sv:56:5
												wire [NUM_OUTPUTS - 1:0] rsp_valid_in;
												// Trace: src/VX_mem_switch.sv:57:5
												wire [(NUM_OUTPUTS * 35) - 1:0] rsp_data_in;
												// Trace: src/VX_mem_switch.sv:58:5
												wire [NUM_OUTPUTS - 1:0] rsp_ready_in;
												// Trace: src/VX_mem_switch.sv:59:5
												wire [0:0] rsp_valid_out;
												// Trace: src/VX_mem_switch.sv:60:5
												wire [34:0] rsp_data_out;
												// Trace: src/VX_mem_switch.sv:61:5
												wire [0:0] rsp_ready_out;
												// Trace: src/VX_mem_switch.sv:62:5
												genvar _gv_i_111;
												for (_gv_i_111 = 0; _gv_i_111 < NUM_OUTPUTS; _gv_i_111 = _gv_i_111 + 1) begin : g_rsp_data_in
													localparam i = _gv_i_111;
													// Trace: src/VX_mem_switch.sv:63:9
													assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_valid;
													// Trace: src/VX_mem_switch.sv:64:9
													assign rsp_data_in[i * 35+:35] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_data;
													// Trace: src/VX_mem_switch.sv:65:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
												end
												// Trace: src/VX_mem_switch.sv:67:5
												VX_stream_arb #(
													.NUM_INPUTS(NUM_OUTPUTS),
													.NUM_OUTPUTS(NUM_INPUTS),
													.DATAW(RSP_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(RSP_OUT_BUF)
												) rsp_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(rsp_valid_in),
													.data_in(rsp_data_in),
													.ready_in(rsp_ready_in),
													.valid_out(rsp_valid_out),
													.data_out(rsp_data_out),
													.ready_out(rsp_ready_out),
													.sel_out()
												);
												// Trace: src/VX_mem_switch.sv:84:5
												genvar _gv_i_112;
												for (_gv_i_112 = 0; _gv_i_112 < NUM_INPUTS; _gv_i_112 = _gv_i_112 + 1) begin : g_rsp_data_out
													localparam i = _gv_i_112;
													// Trace: src/VX_mem_switch.sv:85:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
													// Trace: src/VX_mem_switch.sv:86:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 35+:35];
													// Trace: src/VX_mem_switch.sv:87:9
													assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_bus_in_if].rsp_ready;
												end
											end
											assign core_bus_nc_switch.clk = clk;
											assign core_bus_nc_switch.reset = reset;
											assign core_bus_nc_switch.bus_sel = core_req_nc_sel;
											// Trace: src/VX_cache_bypass.sv:58:5
											// expanded interface instance: core_bus_in_nc_if
											localparam _param_C0263_DATA_SIZE = WORD_SIZE;
											localparam _param_C0263_TAG_WIDTH = CORE_TAG_WIDTH;
											genvar _arr_C0263;
											for (_arr_C0263 = 0; _arr_C0263 <= 0; _arr_C0263 = _arr_C0263 + 1) begin : core_bus_in_nc_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_C0263_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_C0263_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 30;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [72:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [34:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache_bypass.sv:62:5
											genvar _gv_i_57;
											for (_gv_i_57 = 0; _gv_i_57 < NUM_REQS; _gv_i_57 = _gv_i_57 + 1) begin : g_core_bus_nc_switch_if
												localparam i = _gv_i_57;
												// Trace: src/VX_cache_bypass.sv:63:9
												assign core_bus_in_nc_if[i].req_valid = core_bus_nc_switch_if[0 + i].req_valid;
												// Trace: src/VX_cache_bypass.sv:64:9
												assign core_bus_in_nc_if[i].req_data = core_bus_nc_switch_if[0 + i].req_data;
												// Trace: src/VX_cache_bypass.sv:65:9
												assign core_bus_nc_switch_if[0 + i].req_ready = core_bus_in_nc_if[i].req_ready;
												// Trace: src/VX_cache_bypass.sv:66:9
												assign core_bus_nc_switch_if[0 + i].rsp_valid = core_bus_in_nc_if[i].rsp_valid;
												// Trace: src/VX_cache_bypass.sv:67:9
												assign core_bus_nc_switch_if[0 + i].rsp_data = core_bus_in_nc_if[i].rsp_data;
												// Trace: src/VX_cache_bypass.sv:68:9
												assign core_bus_in_nc_if[i].rsp_ready = core_bus_nc_switch_if[0 + i].rsp_ready;
												if (CACHE_ENABLE) begin : g_cache
													// Trace: src/VX_cache_bypass.sv:70:13
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = core_bus_nc_switch_if[1 + i].req_valid;
													// Trace: src/VX_cache_bypass.sv:71:13
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = core_bus_nc_switch_if[1 + i].req_data;
													// Trace: src/VX_cache_bypass.sv:72:13
													assign core_bus_nc_switch_if[1 + i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_ready;
													// Trace: src/VX_cache_bypass.sv:73:13
													assign core_bus_nc_switch_if[1 + i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_valid;
													// Trace: src/VX_cache_bypass.sv:74:13
													assign core_bus_nc_switch_if[1 + i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_data;
													// Trace: src/VX_cache_bypass.sv:75:13
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = core_bus_nc_switch_if[1 + i].rsp_ready;
												end
												else begin : g_no_cache
													// Trace: src/VX_cache_bypass.sv:77:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = 0;
													// Trace: src/VX_cache_bypass.sv:78:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = 1'sb0;
													// Trace: src/VX_cache_bypass.sv:79:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = 0;
												end
											end
											// Trace: src/VX_cache_bypass.sv:82:5
											// expanded interface instance: core_bus_nc_arb_if
											localparam _param_D50AC_DATA_SIZE = WORD_SIZE;
											localparam _param_D50AC_TAG_WIDTH = MEM_TAG_NC1_WIDTH;
											genvar _arr_D50AC;
											for (_arr_D50AC = 0; _arr_D50AC <= 0; _arr_D50AC = _arr_D50AC + 1) begin : core_bus_nc_arb_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_D50AC_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_D50AC_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 30;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [72:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [34:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache_bypass.sv:86:5
											// expanded module instance: core_bus_nc_arb
											localparam _bbase_1376F_bus_in_if = 0;
											localparam _bbase_1376F_bus_out_if = 0;
											localparam _param_1376F_NUM_INPUTS = NUM_REQS;
											localparam _param_1376F_NUM_OUTPUTS = MEM_PORTS;
											localparam _param_1376F_DATA_SIZE = WORD_SIZE;
											localparam _param_1376F_TAG_WIDTH = CORE_TAG_WIDTH;
											localparam _param_1376F_TAG_SEL_IDX = TAG_SEL_IDX;
											localparam _param_1376F_ARBITER = (CACHE_ENABLE ? "P" : "R");
											localparam _param_1376F_REQ_OUT_BUF = 0;
											localparam _param_1376F_RSP_OUT_BUF = 0;
											if (1) begin : core_bus_nc_arb
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_arb.sv:2:15
												localparam NUM_INPUTS = _param_1376F_NUM_INPUTS;
												// Trace: src/VX_mem_arb.sv:3:15
												localparam NUM_OUTPUTS = _param_1376F_NUM_OUTPUTS;
												// Trace: src/VX_mem_arb.sv:4:15
												localparam DATA_SIZE = _param_1376F_DATA_SIZE;
												// Trace: src/VX_mem_arb.sv:5:15
												localparam TAG_WIDTH = _param_1376F_TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:6:15
												localparam TAG_SEL_IDX = _param_1376F_TAG_SEL_IDX;
												// Trace: src/VX_mem_arb.sv:7:15
												localparam REQ_OUT_BUF = _param_1376F_REQ_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:8:15
												localparam RSP_OUT_BUF = _param_1376F_RSP_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:9:15
												localparam ARBITER = _param_1376F_ARBITER;
												// Trace: src/VX_mem_arb.sv:10:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_arb.sv:11:15
												localparam ADDR_WIDTH = 30;
												// Trace: src/VX_mem_arb.sv:12:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_arb.sv:14:5
												wire clk;
												// Trace: src/VX_mem_arb.sv:15:5
												wire reset;
												// Trace: src/VX_mem_arb.sv:16:5
												localparam _mbase_bus_in_if = 0;
												// Trace: src/VX_mem_arb.sv:17:5
												localparam _mbase_bus_out_if = 0;
												// Trace: src/VX_mem_arb.sv:19:5
												localparam DATA_WIDTH = 32;
												// Trace: src/VX_mem_arb.sv:20:5
												localparam LOG_NUM_REQS = 0;
												// Trace: src/VX_mem_arb.sv:21:5
												localparam REQ_DATAW = 73;
												// Trace: src/VX_mem_arb.sv:22:5
												localparam RSP_DATAW = 35;
												// Trace: src/VX_mem_arb.sv:23:5
												localparam SEL_COUNT = NUM_OUTPUTS;
												// Trace: src/VX_mem_arb.sv:24:5
												wire [0:0] req_valid_in;
												// Trace: src/VX_mem_arb.sv:25:5
												wire [72:0] req_data_in;
												// Trace: src/VX_mem_arb.sv:26:5
												wire [0:0] req_ready_in;
												// Trace: src/VX_mem_arb.sv:27:5
												wire [0:0] req_valid_out;
												// Trace: src/VX_mem_arb.sv:28:5
												wire [72:0] req_data_out;
												// Trace: src/VX_mem_arb.sv:29:5
												wire [0:0] req_sel_out;
												// Trace: src/VX_mem_arb.sv:30:5
												wire [0:0] req_ready_out;
												// Trace: src/VX_mem_arb.sv:31:5
												genvar _gv_i_183;
												for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
													localparam i = _gv_i_183;
													// Trace: src/VX_mem_arb.sv:32:9
													assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_valid;
													// Trace: src/VX_mem_arb.sv:33:9
													assign req_data_in[i * 73+:73] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_data;
													// Trace: src/VX_mem_arb.sv:34:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
												end
												// Trace: src/VX_mem_arb.sv:36:5
												VX_stream_arb #(
													.NUM_INPUTS(NUM_INPUTS),
													.NUM_OUTPUTS(NUM_OUTPUTS),
													.DATAW(REQ_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(REQ_OUT_BUF)
												) req_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(req_valid_in),
													.ready_in(req_ready_in),
													.data_in(req_data_in),
													.data_out(req_data_out),
													.sel_out(req_sel_out),
													.valid_out(req_valid_out),
													.ready_out(req_ready_out)
												);
												// Trace: src/VX_mem_arb.sv:53:5
												genvar _gv_i_184;
												for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
													localparam i = _gv_i_184;
													// Trace: src/VX_mem_arb.sv:54:9
													wire [2:0] req_tag_out;
													// Trace: src/VX_mem_arb.sv:55:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
													// Trace: src/VX_mem_arb.sv:56:9
													assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[72], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[71-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[41-:32], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[9-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[5-:3], req_tag_out} = req_data_out[i * 73+:73];
													// Trace: src/VX_mem_arb.sv:64:9
													assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_ready;
													if (1) begin : g_req_tag_out
														// Trace: src/VX_mem_arb.sv:76:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[2-:3] = req_tag_out;
													end
												end
												// Trace: src/VX_mem_arb.sv:79:5
												wire [0:0] rsp_valid_out;
												// Trace: src/VX_mem_arb.sv:80:5
												wire [34:0] rsp_data_out;
												// Trace: src/VX_mem_arb.sv:81:5
												wire [0:0] rsp_ready_out;
												// Trace: src/VX_mem_arb.sv:82:5
												wire [0:0] rsp_valid_in;
												// Trace: src/VX_mem_arb.sv:83:5
												wire [34:0] rsp_data_in;
												// Trace: src/VX_mem_arb.sv:84:5
												wire [0:0] rsp_ready_in;
												// Trace: src/VX_mem_arb.sv:85:5
												if (1) begin : g_rsp_arb
													genvar _gv_i_186;
													for (_gv_i_186 = 0; _gv_i_186 < NUM_OUTPUTS; _gv_i_186 = _gv_i_186 + 1) begin : g_rsp_data_in
														localparam i = _gv_i_186;
														// Trace: src/VX_mem_arb.sv:120:13
														assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_valid;
														// Trace: src/VX_mem_arb.sv:121:13
														assign rsp_data_in[i * 35+:35] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_data;
														// Trace: src/VX_mem_arb.sv:122:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
													end
													// Trace: src/VX_mem_arb.sv:124:9
													VX_stream_arb #(
														.NUM_INPUTS(NUM_OUTPUTS),
														.NUM_OUTPUTS(NUM_INPUTS),
														.DATAW(RSP_DATAW),
														.ARBITER(ARBITER),
														.OUT_BUF(RSP_OUT_BUF)
													) req_arb(
														.clk(clk),
														.reset(reset),
														.valid_in(rsp_valid_in),
														.ready_in(rsp_ready_in),
														.data_in(rsp_data_in),
														.data_out(rsp_data_out),
														.valid_out(rsp_valid_out),
														.ready_out(rsp_ready_out),
														.sel_out()
													);
												end
												// Trace: src/VX_mem_arb.sv:142:5
												genvar _gv_i_187;
												for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
													localparam i = _gv_i_187;
													// Trace: src/VX_mem_arb.sv:143:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
													// Trace: src/VX_mem_arb.sv:144:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 35+:35];
													// Trace: src/VX_mem_arb.sv:145:9
													assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_ready;
												end
											end
											assign core_bus_nc_arb.clk = clk;
											assign core_bus_nc_arb.reset = reset;
											// Trace: src/VX_cache_bypass.sv:101:5
											// expanded interface instance: mem_bus_out_nc_if
											localparam _param_0061C_DATA_SIZE = LINE_SIZE;
											localparam _param_0061C_TAG_WIDTH = MEM_TAG_NC2_WIDTH;
											genvar _arr_0061C;
											for (_arr_0061C = 0; _arr_0061C <= 0; _arr_0061C = _arr_0061C + 1) begin : mem_bus_out_nc_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_0061C_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_0061C_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [612:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [518:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache_bypass.sv:105:5
											genvar _gv_i_58;
											localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
											localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
											for (_gv_i_58 = 0; _gv_i_58 < MEM_PORTS; _gv_i_58 = _gv_i_58 + 1) begin : g_mem_bus_out_nc
												localparam i = _gv_i_58;
												// Trace: src/VX_cache_bypass.sv:106:9
												wire core_req_nc_arb_rw;
												// Trace: src/VX_cache_bypass.sv:107:9
												wire [3:0] core_req_nc_arb_byteen;
												// Trace: src/VX_cache_bypass.sv:108:9
												wire [29:0] core_req_nc_arb_addr;
												// Trace: src/VX_cache_bypass.sv:109:9
												wire [2:0] core_req_nc_arb_flags;
												// Trace: src/VX_cache_bypass.sv:110:9
												wire [31:0] core_req_nc_arb_data;
												// Trace: src/VX_cache_bypass.sv:111:9
												wire [2:0] core_req_nc_arb_tag;
												// Trace: src/VX_cache_bypass.sv:112:9
												assign {core_req_nc_arb_rw, core_req_nc_arb_addr, core_req_nc_arb_data, core_req_nc_arb_byteen, core_req_nc_arb_flags, core_req_nc_arb_tag} = core_bus_nc_arb_if[i].req_data;
												// Trace: src/VX_cache_bypass.sv:120:9
												wire [25:0] core_req_nc_arb_addr_w;
												// Trace: src/VX_cache_bypass.sv:121:9
												reg [63:0] core_req_nc_arb_byteen_w;
												// Trace: src/VX_cache_bypass.sv:122:9
												reg [511:0] core_req_nc_arb_data_w;
												// Trace: src/VX_cache_bypass.sv:123:9
												wire [31:0] core_rsp_nc_arb_data_w;
												// Trace: src/VX_cache_bypass.sv:124:9
												wire [6:0] core_req_nc_arb_tag_w;
												// Trace: src/VX_cache_bypass.sv:125:9
												wire [2:0] core_rsp_nc_arb_tag_w;
												if (1) begin : g_multi_word_line
													// Trace: src/VX_cache_bypass.sv:127:13
													wire [3:0] rsp_wsel;
													// Trace: src/VX_cache_bypass.sv:128:13
													wire [3:0] req_wsel = core_req_nc_arb_addr[3:0];
													// Trace: src/VX_cache_bypass.sv:129:13
													always @(*) begin
														// Trace: src/VX_cache_bypass.sv:130:17
														core_req_nc_arb_byteen_w = 1'sb0;
														// Trace: src/VX_cache_bypass.sv:131:17
														core_req_nc_arb_byteen_w[req_wsel * 4+:4] = core_req_nc_arb_byteen;
														// Trace: src/VX_cache_bypass.sv:132:17
														core_req_nc_arb_data_w = 1'sbx;
														// Trace: src/VX_cache_bypass.sv:133:17
														core_req_nc_arb_data_w[req_wsel * 32+:32] = core_req_nc_arb_data;
													end
													// Trace: src/VX_cache_bypass.sv:135:13
													VX_bits_insert #(
														.N(MEM_TAG_NC1_WIDTH),
														.S(WSEL_BITS),
														.POS(TAG_SEL_IDX)
													) wsel_insert(
														.data_in(core_req_nc_arb_tag),
														.ins_in(req_wsel),
														.data_out(core_req_nc_arb_tag_w)
													);
													// Trace: src/VX_cache_bypass.sv:144:13
													VX_bits_remove #(
														.N(MEM_TAG_NC2_WIDTH),
														.S(WSEL_BITS),
														.POS(TAG_SEL_IDX)
													) wsel_remove(
														.data_in(mem_bus_out_nc_if[i].rsp_data[6-:7]),
														.sel_out(rsp_wsel),
														.data_out(core_rsp_nc_arb_tag_w)
													);
													// Trace: src/VX_cache_bypass.sv:153:13
													assign core_req_nc_arb_addr_w = core_req_nc_arb_addr[WSEL_BITS+:MEM_ADDR_WIDTH];
													// Trace: src/VX_cache_bypass.sv:154:13
													assign core_rsp_nc_arb_data_w = mem_bus_out_nc_if[i].rsp_data[7 + (rsp_wsel * CORE_DATA_WIDTH)+:CORE_DATA_WIDTH];
												end
												// Trace: src/VX_cache_bypass.sv:163:9
												assign mem_bus_out_nc_if[i].req_valid = core_bus_nc_arb_if[i].req_valid;
												// Trace: src/VX_cache_bypass.sv:164:9
												assign mem_bus_out_nc_if[i].req_data = {core_req_nc_arb_rw, core_req_nc_arb_addr_w, core_req_nc_arb_data_w, core_req_nc_arb_byteen_w, core_req_nc_arb_flags, core_req_nc_arb_tag_w};
												// Trace: src/VX_cache_bypass.sv:172:9
												assign core_bus_nc_arb_if[i].req_ready = mem_bus_out_nc_if[i].req_ready;
												// Trace: src/VX_cache_bypass.sv:173:9
												assign core_bus_nc_arb_if[i].rsp_valid = mem_bus_out_nc_if[i].rsp_valid;
												// Trace: src/VX_cache_bypass.sv:174:9
												assign core_bus_nc_arb_if[i].rsp_data = {core_rsp_nc_arb_data_w, core_rsp_nc_arb_tag_w};
												// Trace: src/VX_cache_bypass.sv:178:9
												assign mem_bus_out_nc_if[i].rsp_ready = core_bus_nc_arb_if[i].rsp_ready;
											end
											// Trace: src/VX_cache_bypass.sv:180:5
											// expanded interface instance: mem_bus_out_src_if
											localparam _param_913F6_DATA_SIZE = LINE_SIZE;
											localparam _param_913F6_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
											genvar _arr_913F6;
											for (_arr_913F6 = 0; _arr_913F6 <= (((CACHE_ENABLE ? 2 : 1) * MEM_PORTS) - 1); _arr_913F6 = _arr_913F6 + 1) begin : mem_bus_out_src_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_913F6_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_913F6_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [612:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [518:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache_bypass.sv:184:5
											genvar _gv_i_59;
											for (_gv_i_59 = 0; _gv_i_59 < MEM_PORTS; _gv_i_59 = _gv_i_59 + 1) begin : g_mem_bus_out_src
												localparam i = _gv_i_59;
												// Trace: src/VX_cache_bypass.sv:186:5
												assign mem_bus_out_src_if[0 + i].req_valid = mem_bus_out_nc_if[i].req_valid;
												// Trace: src/VX_cache_bypass.sv:187:5
												assign mem_bus_out_src_if[0 + i].req_data[612] = mem_bus_out_nc_if[i].req_data[612];
												// Trace: src/VX_cache_bypass.sv:188:5
												assign mem_bus_out_src_if[0 + i].req_data[611-:26] = mem_bus_out_nc_if[i].req_data[611-:26];
												// Trace: src/VX_cache_bypass.sv:189:5
												assign mem_bus_out_src_if[0 + i].req_data[585-:512] = mem_bus_out_nc_if[i].req_data[585-:512];
												// Trace: src/VX_cache_bypass.sv:190:5
												assign mem_bus_out_src_if[0 + i].req_data[73-:64] = mem_bus_out_nc_if[i].req_data[73-:64];
												// Trace: src/VX_cache_bypass.sv:191:5
												assign mem_bus_out_src_if[0 + i].req_data[9-:3] = mem_bus_out_nc_if[i].req_data[9-:3];
												if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk1
													if (1) begin : genblk1
														if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
															// Trace: src/VX_cache_bypass.sv:195:17
															assign mem_bus_out_src_if[0 + i].req_data[6-:7] = {mem_bus_out_nc_if[i].req_data[6-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_NC2_WIDTH {1'b0}}, mem_bus_out_nc_if[i].req_data[5-:6]};
														end
														else begin : genblk1
															// Trace: src/VX_cache_bypass.sv:197:17
															assign mem_bus_out_src_if[0 + i].req_data[6-:7] = {mem_bus_out_nc_if[i].req_data[6-:1], mem_bus_out_nc_if[i].req_data[(MEM_TAG_OUT_WIDTH - VX_gpu_pkg_UUID_WIDTH) - 1:0]};
														end
													end
												end
												else begin : genblk1
													// Trace: src/VX_cache_bypass.sv:207:9
													assign mem_bus_out_src_if[0 + i].req_data[6-:7] = mem_bus_out_nc_if[i].req_data[6-:7];
												end
												// Trace: src/VX_cache_bypass.sv:209:5
												assign mem_bus_out_nc_if[i].req_ready = mem_bus_out_src_if[0 + i].req_ready;
												// Trace: src/VX_cache_bypass.sv:210:5
												assign mem_bus_out_nc_if[i].rsp_valid = mem_bus_out_src_if[0 + i].rsp_valid;
												// Trace: src/VX_cache_bypass.sv:211:5
												assign mem_bus_out_nc_if[i].rsp_data[518-:512] = mem_bus_out_src_if[0 + i].rsp_data[518-:512];
												if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk2
													if (1) begin : genblk1
														if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
															// Trace: src/VX_cache_bypass.sv:215:17
															assign mem_bus_out_nc_if[i].rsp_data[6-:7] = {mem_bus_out_src_if[0 + i].rsp_data[6-:1], mem_bus_out_src_if[0 + i].rsp_data[5:0]};
														end
														else begin : genblk1
															// Trace: src/VX_cache_bypass.sv:217:17
															assign mem_bus_out_nc_if[i].rsp_data[6-:7] = {mem_bus_out_src_if[0 + i].rsp_data[6-:1], {MEM_TAG_NC2_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[0 + i].rsp_data[5-:6]};
														end
													end
												end
												else begin : genblk2
													// Trace: src/VX_cache_bypass.sv:227:9
													assign mem_bus_out_nc_if[i].rsp_data[6-:7] = mem_bus_out_src_if[0 + i].rsp_data[6-:7];
												end
												// Trace: src/VX_cache_bypass.sv:229:5
												assign mem_bus_out_src_if[0 + i].rsp_ready = mem_bus_out_nc_if[i].rsp_ready;
												if (CACHE_ENABLE) begin : g_cache
													// Trace: src/VX_cache_bypass.sv:233:5
													assign mem_bus_out_src_if[1 + i].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_valid;
													// Trace: src/VX_cache_bypass.sv:234:5
													assign mem_bus_out_src_if[1 + i].req_data[612] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[610];
													// Trace: src/VX_cache_bypass.sv:235:5
													assign mem_bus_out_src_if[1 + i].req_data[611-:26] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[609-:26];
													// Trace: src/VX_cache_bypass.sv:236:5
													assign mem_bus_out_src_if[1 + i].req_data[585-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[583-:512];
													// Trace: src/VX_cache_bypass.sv:237:5
													assign mem_bus_out_src_if[1 + i].req_data[73-:64] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[71-:64];
													// Trace: src/VX_cache_bypass.sv:238:5
													assign mem_bus_out_src_if[1 + i].req_data[9-:3] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[7-:3];
													if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk1
														if (1) begin : genblk1
															if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
																// Trace: src/VX_cache_bypass.sv:242:17
																assign mem_bus_out_src_if[1 + i].req_data[6-:7] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_IN_WIDTH {1'b0}}, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[3-:4]};
															end
															else begin : genblk1
																// Trace: src/VX_cache_bypass.sv:244:17
																assign mem_bus_out_src_if[1 + i].req_data[6-:7] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[(MEM_TAG_OUT_WIDTH - VX_gpu_pkg_UUID_WIDTH) - 1:0]};
															end
														end
													end
													else begin : genblk1
														// Trace: src/VX_cache_bypass.sv:254:9
														assign mem_bus_out_src_if[1 + i].req_data[6-:7] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:5];
													end
													// Trace: src/VX_cache_bypass.sv:256:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = mem_bus_out_src_if[1 + i].req_ready;
													// Trace: src/VX_cache_bypass.sv:257:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = mem_bus_out_src_if[1 + i].rsp_valid;
													// Trace: src/VX_cache_bypass.sv:258:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[516-:512] = mem_bus_out_src_if[1 + i].rsp_data[518-:512];
													if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk2
														if (1) begin : genblk1
															if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
																// Trace: src/VX_cache_bypass.sv:262:17
																assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[6-:1], mem_bus_out_src_if[1 + i].rsp_data[3:0]};
															end
															else begin : genblk1
																// Trace: src/VX_cache_bypass.sv:264:17
																assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[6-:1], {MEM_TAG_IN_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[1 + i].rsp_data[5-:6]};
															end
														end
													end
													else begin : genblk2
														// Trace: src/VX_cache_bypass.sv:274:9
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = mem_bus_out_src_if[1 + i].rsp_data[6-:7];
													end
													// Trace: src/VX_cache_bypass.sv:276:5
													assign mem_bus_out_src_if[1 + i].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_ready;
												end
												else begin : g_no_cache
													// Trace: src/VX_cache_bypass.sv:279:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = 0;
													// Trace: src/VX_cache_bypass.sv:280:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = 0;
													// Trace: src/VX_cache_bypass.sv:281:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data = 1'sb0;
												end
											end
											// Trace: src/VX_cache_bypass.sv:284:5
											// expanded module instance: mem_bus_out_arb
											localparam _bbase_B06D0_bus_in_if = 0;
											localparam _bbase_B06D0_bus_out_if = 0;
											localparam _param_B06D0_NUM_INPUTS = (CACHE_ENABLE ? 2 : 1) * MEM_PORTS;
											localparam _param_B06D0_NUM_OUTPUTS = MEM_PORTS;
											localparam _param_B06D0_DATA_SIZE = LINE_SIZE;
											localparam _param_B06D0_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
											localparam _param_B06D0_ARBITER = "R";
											localparam _param_B06D0_REQ_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
											localparam _param_B06D0_RSP_OUT_BUF = 0;
											if (1) begin : mem_bus_out_arb
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_arb.sv:2:15
												localparam NUM_INPUTS = _param_B06D0_NUM_INPUTS;
												// Trace: src/VX_mem_arb.sv:3:15
												localparam NUM_OUTPUTS = _param_B06D0_NUM_OUTPUTS;
												// Trace: src/VX_mem_arb.sv:4:15
												localparam DATA_SIZE = _param_B06D0_DATA_SIZE;
												// Trace: src/VX_mem_arb.sv:5:15
												localparam TAG_WIDTH = _param_B06D0_TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:6:15
												localparam TAG_SEL_IDX = 0;
												// Trace: src/VX_mem_arb.sv:7:15
												localparam REQ_OUT_BUF = _param_B06D0_REQ_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:8:15
												localparam RSP_OUT_BUF = _param_B06D0_RSP_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:9:15
												localparam ARBITER = _param_B06D0_ARBITER;
												// Trace: src/VX_mem_arb.sv:10:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_arb.sv:11:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_arb.sv:12:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_arb.sv:14:5
												wire clk;
												// Trace: src/VX_mem_arb.sv:15:5
												wire reset;
												// Trace: src/VX_mem_arb.sv:16:5
												localparam _mbase_bus_in_if = 0;
												// Trace: src/VX_mem_arb.sv:17:5
												localparam _mbase_bus_out_if = 0;
												// Trace: src/VX_mem_arb.sv:19:5
												localparam DATA_WIDTH = 512;
												// Trace: src/VX_mem_arb.sv:20:5
												localparam LOG_NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? $clog2((NUM_INPUTS + 0) / 1) : 0);
												// Trace: src/VX_mem_arb.sv:21:5
												localparam REQ_DATAW = 606 + TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:22:5
												localparam RSP_DATAW = DATA_WIDTH + TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:23:5
												localparam SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
												// Trace: src/VX_mem_arb.sv:24:5
												wire [NUM_INPUTS - 1:0] req_valid_in;
												// Trace: src/VX_mem_arb.sv:25:5
												wire [(NUM_INPUTS * REQ_DATAW) - 1:0] req_data_in;
												// Trace: src/VX_mem_arb.sv:26:5
												wire [NUM_INPUTS - 1:0] req_ready_in;
												// Trace: src/VX_mem_arb.sv:27:5
												wire [0:0] req_valid_out;
												// Trace: src/VX_mem_arb.sv:28:5
												wire [REQ_DATAW - 1:0] req_data_out;
												// Trace: src/VX_mem_arb.sv:29:5
												wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] req_sel_out;
												// Trace: src/VX_mem_arb.sv:30:5
												wire [0:0] req_ready_out;
												// Trace: src/VX_mem_arb.sv:31:5
												genvar _gv_i_183;
												for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
													localparam i = _gv_i_183;
													// Trace: src/VX_mem_arb.sv:32:9
													assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_valid;
													// Trace: src/VX_mem_arb.sv:33:9
													assign req_data_in[i * 613+:613] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_data;
													// Trace: src/VX_mem_arb.sv:34:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
												end
												// Trace: src/VX_mem_arb.sv:36:5
												VX_stream_arb #(
													.NUM_INPUTS(NUM_INPUTS),
													.NUM_OUTPUTS(NUM_OUTPUTS),
													.DATAW(REQ_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(REQ_OUT_BUF)
												) req_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(req_valid_in),
													.ready_in(req_ready_in),
													.data_in(req_data_in),
													.data_out(req_data_out),
													.sel_out(req_sel_out),
													.valid_out(req_valid_out),
													.ready_out(req_ready_out)
												);
												// Trace: src/VX_mem_arb.sv:53:5
												genvar _gv_i_184;
												for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
													localparam i = _gv_i_184;
													// Trace: src/VX_mem_arb.sv:54:9
													wire [TAG_WIDTH - 1:0] req_tag_out;
													// Trace: src/VX_mem_arb.sv:55:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
													// Trace: src/VX_mem_arb.sv:56:9
													assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[610], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[609-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[583-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[71-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[7-:3], req_tag_out} = req_data_out[i * 613+:613];
													// Trace: src/VX_mem_arb.sv:64:9
													assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
													if (NUM_INPUTS > NUM_OUTPUTS) begin : g_req_tag_sel_out
														// Trace: src/VX_mem_arb.sv:66:13
														VX_bits_insert #(
															.N(TAG_WIDTH),
															.S(LOG_NUM_REQS),
															.POS(TAG_SEL_IDX)
														) bits_insert(
															.data_in(req_tag_out),
															.ins_in(req_sel_out[i * 1+:1]),
															.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[4-:5])
														);
													end
													else begin : g_req_tag_out
														// Trace: src/VX_mem_arb.sv:76:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[4-:5] = req_tag_out;
													end
												end
												// Trace: src/VX_mem_arb.sv:79:5
												wire [NUM_INPUTS - 1:0] rsp_valid_out;
												// Trace: src/VX_mem_arb.sv:80:5
												wire [(NUM_INPUTS * RSP_DATAW) - 1:0] rsp_data_out;
												// Trace: src/VX_mem_arb.sv:81:5
												wire [NUM_INPUTS - 1:0] rsp_ready_out;
												// Trace: src/VX_mem_arb.sv:82:5
												wire [0:0] rsp_valid_in;
												// Trace: src/VX_mem_arb.sv:83:5
												wire [RSP_DATAW - 1:0] rsp_data_in;
												// Trace: src/VX_mem_arb.sv:84:5
												wire [0:0] rsp_ready_in;
												// Trace: src/VX_mem_arb.sv:85:5
												if (NUM_INPUTS > NUM_OUTPUTS) begin : g_rsp_select
													// Trace: src/VX_mem_arb.sv:86:9
													wire [LOG_NUM_REQS - 1:0] rsp_sel_in;
													genvar _gv_i_185;
													for (_gv_i_185 = 0; _gv_i_185 < NUM_OUTPUTS; _gv_i_185 = _gv_i_185 + 1) begin : g_rsp_data_in
														localparam i = _gv_i_185;
														// Trace: src/VX_mem_arb.sv:88:13
														wire [TAG_WIDTH - 1:0] rsp_tag_out;
														// Trace: src/VX_mem_arb.sv:89:13
														VX_bits_remove #(
															.N(TAG_WIDTH + LOG_NUM_REQS),
															.S(LOG_NUM_REQS),
															.POS(TAG_SEL_IDX)
														) bits_remove(
															.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[4-:5]),
															.sel_out(rsp_sel_in[i * 1+:1]),
															.data_out(rsp_tag_out)
														);
														// Trace: src/VX_mem_arb.sv:98:13
														assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
														// Trace: src/VX_mem_arb.sv:99:13
														assign rsp_data_in[i * 519+:519] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[516-:512], rsp_tag_out};
														// Trace: src/VX_mem_arb.sv:100:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
													end
													// Trace: src/VX_mem_arb.sv:102:9
													VX_stream_switch #(
														.NUM_INPUTS(NUM_OUTPUTS),
														.NUM_OUTPUTS(NUM_INPUTS),
														.DATAW(RSP_DATAW),
														.OUT_BUF(RSP_OUT_BUF)
													) rsp_switch(
														.clk(clk),
														.reset(reset),
														.sel_in(rsp_sel_in),
														.valid_in(rsp_valid_in),
														.ready_in(rsp_ready_in),
														.data_in(rsp_data_in),
														.data_out(rsp_data_out),
														.valid_out(rsp_valid_out),
														.ready_out(rsp_ready_out)
													);
												end
												else begin : g_rsp_arb
													genvar _gv_i_186;
													for (_gv_i_186 = 0; _gv_i_186 < NUM_OUTPUTS; _gv_i_186 = _gv_i_186 + 1) begin : g_rsp_data_in
														localparam i = _gv_i_186;
														// Trace: src/VX_mem_arb.sv:120:13
														assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
														// Trace: src/VX_mem_arb.sv:121:13
														assign rsp_data_in[i * 519+:519] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
														// Trace: src/VX_mem_arb.sv:122:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
													end
													// Trace: src/VX_mem_arb.sv:124:9
													VX_stream_arb #(
														.NUM_INPUTS(NUM_OUTPUTS),
														.NUM_OUTPUTS(NUM_INPUTS),
														.DATAW(RSP_DATAW),
														.ARBITER(ARBITER),
														.OUT_BUF(RSP_OUT_BUF)
													) req_arb(
														.clk(clk),
														.reset(reset),
														.valid_in(rsp_valid_in),
														.ready_in(rsp_ready_in),
														.data_in(rsp_data_in),
														.data_out(rsp_data_out),
														.valid_out(rsp_valid_out),
														.ready_out(rsp_ready_out),
														.sel_out()
													);
												end
												// Trace: src/VX_mem_arb.sv:142:5
												genvar _gv_i_187;
												for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
													localparam i = _gv_i_187;
													// Trace: src/VX_mem_arb.sv:143:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
													// Trace: src/VX_mem_arb.sv:144:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 519+:519];
													// Trace: src/VX_mem_arb.sv:145:9
													assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_ready;
												end
											end
											assign mem_bus_out_arb.clk = clk;
											assign mem_bus_out_arb.reset = reset;
										end
										assign cache_bypass.clk = clk;
										assign cache_bypass.reset = reset;
									end
									else begin : g_no_bypass
										genvar _gv_i_38;
										for (_gv_i_38 = 0; _gv_i_38 < NUM_REQS; _gv_i_38 = _gv_i_38 + 1) begin : g_core_bus_cache_if
											localparam i = _gv_i_38;
											// Trace: src/VX_cache_wrap.sv:73:5
											assign core_bus_cache_if[i].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_if].req_valid;
											// Trace: src/VX_cache_wrap.sv:74:5
											assign core_bus_cache_if[i].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_if].req_data;
											// Trace: src/VX_cache_wrap.sv:75:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_if].req_ready = core_bus_cache_if[i].req_ready;
											// Trace: src/VX_cache_wrap.sv:76:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_if].rsp_valid = core_bus_cache_if[i].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:77:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_if].rsp_data = core_bus_cache_if[i].rsp_data;
											// Trace: src/VX_cache_wrap.sv:78:5
											assign core_bus_cache_if[i].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.arb_core_bus_if[i + _mbase_core_bus_if].rsp_ready;
										end
										genvar _gv_i_39;
										for (_gv_i_39 = 0; _gv_i_39 < MEM_PORTS; _gv_i_39 = _gv_i_39 + 1) begin : g_mem_bus_tmp_if
											localparam i = _gv_i_39;
											// Trace: src/VX_cache_wrap.sv:81:5
											assign mem_bus_tmp_if[i].req_valid = mem_bus_cache_if[i].req_valid;
											// Trace: src/VX_cache_wrap.sv:82:5
											assign mem_bus_tmp_if[i].req_data = mem_bus_cache_if[i].req_data;
											// Trace: src/VX_cache_wrap.sv:83:5
											assign mem_bus_cache_if[i].req_ready = mem_bus_tmp_if[i].req_ready;
											// Trace: src/VX_cache_wrap.sv:84:5
											assign mem_bus_cache_if[i].rsp_valid = mem_bus_tmp_if[i].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:85:5
											assign mem_bus_cache_if[i].rsp_data = mem_bus_tmp_if[i].rsp_data;
											// Trace: src/VX_cache_wrap.sv:86:5
											assign mem_bus_tmp_if[i].rsp_ready = mem_bus_cache_if[i].rsp_ready;
										end
									end
									// Trace: src/VX_cache_wrap.sv:89:5
									genvar _gv_i_40;
									for (_gv_i_40 = 0; _gv_i_40 < MEM_PORTS; _gv_i_40 = _gv_i_40 + 1) begin : g_mem_bus_if
										localparam i = _gv_i_40;
										if (WRITE_ENABLE) begin : g_we
											// Trace: src/VX_cache_wrap.sv:91:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
											// Trace: src/VX_cache_wrap.sv:92:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[i].req_data;
											// Trace: src/VX_cache_wrap.sv:93:5
											assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
											// Trace: src/VX_cache_wrap.sv:94:5
											assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:95:5
											assign mem_bus_tmp_if[i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
											// Trace: src/VX_cache_wrap.sv:96:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
										end
										else begin : g_ro
											// Trace: src/VX_cache_wrap.sv:98:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
											// Trace: src/VX_cache_wrap.sv:99:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[610] = 0;
											// Trace: src/VX_cache_wrap.sv:100:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[609-:26] = mem_bus_tmp_if[i].req_data[609-:26];
											// Trace: src/VX_cache_wrap.sv:101:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[583-:512] = 1'sb0;
											// Trace: src/VX_cache_wrap.sv:102:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[71-:64] = 1'sb1;
											// Trace: src/VX_cache_wrap.sv:103:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[7-:3] = mem_bus_tmp_if[i].req_data[7-:3];
											// Trace: src/VX_cache_wrap.sv:104:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[4-:5] = mem_bus_tmp_if[i].req_data[4-:5];
											// Trace: src/VX_cache_wrap.sv:105:5
											assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
											// Trace: src/VX_cache_wrap.sv:106:5
											assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:107:5
											assign mem_bus_tmp_if[i].rsp_data[516-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[516-:512];
											// Trace: src/VX_cache_wrap.sv:108:5
											assign mem_bus_tmp_if[i].rsp_data[4-:5] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[4-:5];
											// Trace: src/VX_cache_wrap.sv:109:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
										end
									end
									// Trace: src/VX_cache_wrap.sv:112:5
									if (1) begin : g_cache
										// Trace: src/VX_cache_wrap.sv:113:9
										// expanded module instance: cache
										localparam _bbase_90EE2_core_bus_if = 0;
										localparam _bbase_90EE2_mem_bus_if = 0;
										localparam _param_90EE2_INSTANCE_ID = INSTANCE_ID;
										localparam _param_90EE2_CACHE_SIZE = CACHE_SIZE;
										localparam _param_90EE2_LINE_SIZE = LINE_SIZE;
										localparam _param_90EE2_NUM_BANKS = NUM_BANKS;
										localparam _param_90EE2_NUM_WAYS = NUM_WAYS;
										localparam _param_90EE2_WORD_SIZE = WORD_SIZE;
										localparam _param_90EE2_NUM_REQS = NUM_REQS;
										localparam _param_90EE2_MEM_PORTS = MEM_PORTS;
										localparam _param_90EE2_WRITE_ENABLE = WRITE_ENABLE;
										localparam _param_90EE2_WRITEBACK = WRITEBACK;
										localparam _param_90EE2_DIRTY_BYTES = DIRTY_BYTES;
										localparam _param_90EE2_REPL_POLICY = REPL_POLICY;
										localparam _param_90EE2_CRSQ_SIZE = CRSQ_SIZE;
										localparam _param_90EE2_MSHR_SIZE = MSHR_SIZE;
										localparam _param_90EE2_MRSQ_SIZE = MRSQ_SIZE;
										localparam _param_90EE2_MREQ_SIZE = MREQ_SIZE;
										localparam _param_90EE2_TAG_WIDTH = TAG_WIDTH;
										localparam _param_90EE2_CORE_OUT_BUF = (BYPASS_ENABLE ? 1 : CORE_OUT_BUF);
										localparam _param_90EE2_MEM_OUT_BUF = (BYPASS_ENABLE ? 1 : MEM_OUT_BUF);
										if (1) begin : cache
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_cache.sv:2:15
											localparam INSTANCE_ID = _param_90EE2_INSTANCE_ID;
											// Trace: src/VX_cache.sv:3:15
											localparam NUM_REQS = _param_90EE2_NUM_REQS;
											// Trace: src/VX_cache.sv:4:15
											localparam MEM_PORTS = _param_90EE2_MEM_PORTS;
											// Trace: src/VX_cache.sv:5:15
											localparam CACHE_SIZE = _param_90EE2_CACHE_SIZE;
											// Trace: src/VX_cache.sv:6:15
											localparam LINE_SIZE = _param_90EE2_LINE_SIZE;
											// Trace: src/VX_cache.sv:7:15
											localparam NUM_BANKS = _param_90EE2_NUM_BANKS;
											// Trace: src/VX_cache.sv:8:15
											localparam NUM_WAYS = _param_90EE2_NUM_WAYS;
											// Trace: src/VX_cache.sv:9:15
											localparam WORD_SIZE = _param_90EE2_WORD_SIZE;
											// Trace: src/VX_cache.sv:10:15
											localparam CRSQ_SIZE = _param_90EE2_CRSQ_SIZE;
											// Trace: src/VX_cache.sv:11:15
											localparam MSHR_SIZE = _param_90EE2_MSHR_SIZE;
											// Trace: src/VX_cache.sv:12:15
											localparam MRSQ_SIZE = _param_90EE2_MRSQ_SIZE;
											// Trace: src/VX_cache.sv:13:15
											localparam MREQ_SIZE = _param_90EE2_MREQ_SIZE;
											// Trace: src/VX_cache.sv:14:15
											localparam WRITE_ENABLE = _param_90EE2_WRITE_ENABLE;
											// Trace: src/VX_cache.sv:15:15
											localparam WRITEBACK = _param_90EE2_WRITEBACK;
											// Trace: src/VX_cache.sv:16:15
											localparam DIRTY_BYTES = _param_90EE2_DIRTY_BYTES;
											// Trace: src/VX_cache.sv:17:15
											localparam REPL_POLICY = _param_90EE2_REPL_POLICY;
											// Trace: src/VX_cache.sv:18:15
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam TAG_WIDTH = _param_90EE2_TAG_WIDTH;
											// Trace: src/VX_cache.sv:19:15
											localparam CORE_OUT_BUF = _param_90EE2_CORE_OUT_BUF;
											// Trace: src/VX_cache.sv:20:15
											localparam MEM_OUT_BUF = _param_90EE2_MEM_OUT_BUF;
											// Trace: src/VX_cache.sv:22:5
											wire clk;
											// Trace: src/VX_cache.sv:23:5
											wire reset;
											// Trace: src/VX_cache.sv:24:5
											localparam _mbase_core_bus_if = 0;
											// Trace: src/VX_cache.sv:25:5
											localparam _mbase_mem_bus_if = 0;
											// Trace: src/VX_cache.sv:27:5
											localparam REQ_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:28:5
											localparam WORD_SEL_WIDTH = 4;
											// Trace: src/VX_cache.sv:29:5
											localparam MSHR_ADDR_WIDTH = 4;
											// Trace: src/VX_cache.sv:30:5
											localparam MEM_TAG_WIDTH = 5;
											// Trace: src/VX_cache.sv:32:5
											localparam WORDS_PER_LINE = 16;
											// Trace: src/VX_cache.sv:33:5
											localparam WORD_WIDTH = 32;
											// Trace: src/VX_cache.sv:34:5
											localparam WORD_SEL_BITS = 4;
											// Trace: src/VX_cache.sv:35:5
											localparam BANK_SEL_BITS = 0;
											// Trace: src/VX_cache.sv:36:5
											localparam BANK_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:37:5
											localparam LINE_ADDR_WIDTH = 26;
											// Trace: src/VX_cache.sv:38:5
											localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
											localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
											localparam CORE_REQ_DATAW = 73;
											// Trace: src/VX_cache.sv:39:5
											localparam CORE_RSP_DATAW = 35;
											// Trace: src/VX_cache.sv:40:5
											localparam BANK_MEM_TAG_WIDTH = 5;
											// Trace: src/VX_cache.sv:41:5
											localparam MEM_REQ_DATAW = 611;
											// Trace: src/VX_cache.sv:42:5
											localparam MEM_RSP_DATAW = 517;
											// Trace: src/VX_cache.sv:43:5
											localparam MEM_PORTS_SEL_BITS = 0;
											// Trace: src/VX_cache.sv:44:5
											localparam MEM_PORTS_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:45:5
											localparam MEM_ARB_SEL_BITS = 0;
											// Trace: src/VX_cache.sv:46:5
											localparam MEM_ARB_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:47:5
											localparam REQ_XBAR_BUF = 0;
											// Trace: src/VX_cache.sv:48:5
											localparam CORE_RSP_BUF_ENABLE = 1'd0;
											// Trace: src/VX_cache.sv:49:5
											localparam MEM_REQ_BUF_ENABLE = 1'd0;
											// Trace: src/VX_cache.sv:50:5
											// expanded interface instance: core_bus2_if
											localparam _param_9260A_DATA_SIZE = WORD_SIZE;
											localparam _param_9260A_TAG_WIDTH = TAG_WIDTH;
											genvar _arr_9260A;
											for (_arr_9260A = 0; _arr_9260A <= 0; _arr_9260A = _arr_9260A + 1) begin : core_bus2_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_9260A_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_9260A_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 30;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [72:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [34:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache.sv:54:5
											wire [0:0] per_bank_flush_begin;
											// Trace: src/VX_cache.sv:55:5
											wire [0:0] flush_uuid;
											// Trace: src/VX_cache.sv:56:5
											wire [0:0] per_bank_flush_end;
											// Trace: src/VX_cache.sv:57:5
											wire [0:0] per_bank_core_req_fire;
											// Trace: src/VX_cache.sv:58:5
											// expanded module instance: cache_init
											localparam _bbase_3B3F2_core_bus_in_if = 0;
											localparam _bbase_3B3F2_core_bus_out_if = 0;
											localparam _param_3B3F2_NUM_REQS = NUM_REQS;
											localparam _param_3B3F2_NUM_BANKS = NUM_BANKS;
											localparam _param_3B3F2_TAG_WIDTH = TAG_WIDTH;
											localparam _param_3B3F2_BANK_SEL_LATENCY = 0;
											if (1) begin : cache_init
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_cache_init.sv:2:15
												localparam NUM_REQS = _param_3B3F2_NUM_REQS;
												// Trace: src/VX_cache_init.sv:3:15
												localparam NUM_BANKS = _param_3B3F2_NUM_BANKS;
												// Trace: src/VX_cache_init.sv:4:15
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam TAG_WIDTH = _param_3B3F2_TAG_WIDTH;
												// Trace: src/VX_cache_init.sv:5:15
												localparam BANK_SEL_LATENCY = _param_3B3F2_BANK_SEL_LATENCY;
												// Trace: src/VX_cache_init.sv:7:5
												wire clk;
												// Trace: src/VX_cache_init.sv:8:5
												wire reset;
												// Trace: src/VX_cache_init.sv:9:5
												localparam _mbase_core_bus_in_if = 0;
												// Trace: src/VX_cache_init.sv:10:5
												localparam _mbase_core_bus_out_if = 0;
												// Trace: src/VX_cache_init.sv:11:5
												wire [0:0] bank_req_fire;
												// Trace: src/VX_cache_init.sv:12:5
												wire [0:0] flush_begin;
												// Trace: src/VX_cache_init.sv:13:5
												wire [0:0] flush_uuid;
												// Trace: src/VX_cache_init.sv:14:5
												wire [0:0] flush_end;
												// Trace: src/VX_cache_init.sv:16:5
												localparam STATE_IDLE = 0;
												// Trace: src/VX_cache_init.sv:17:5
												localparam STATE_WAIT1 = 1;
												// Trace: src/VX_cache_init.sv:18:5
												localparam STATE_FLUSH = 2;
												// Trace: src/VX_cache_init.sv:19:5
												localparam STATE_WAIT2 = 3;
												// Trace: src/VX_cache_init.sv:20:5
												localparam STATE_DONE = 4;
												// Trace: src/VX_cache_init.sv:21:5
												reg [2:0] state;
												reg [2:0] state_n;
												// Trace: src/VX_cache_init.sv:22:5
												wire no_inflight_reqs;
												// Trace: src/VX_cache_init.sv:23:5
												if (1) begin : g_no_bank_sel_latency
													// Trace: src/VX_cache_init.sv:62:9
													assign no_inflight_reqs = 0;
												end
												// Trace: src/VX_cache_init.sv:64:5
												reg [0:0] flush_done;
												reg [0:0] flush_done_n;
												// Trace: src/VX_cache_init.sv:65:5
												wire [0:0] flush_req_mask;
												// Trace: src/VX_cache_init.sv:66:5
												genvar _gv_i_215;
												localparam VX_gpu_pkg_MEM_REQ_FLAG_FLUSH = 0;
												for (_gv_i_215 = 0; _gv_i_215 < NUM_REQS; _gv_i_215 = _gv_i_215 + 1) begin : g_flush_req_mask
													localparam i = _gv_i_215;
													// Trace: src/VX_cache_init.sv:67:9
													assign flush_req_mask[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_data[3];
												end
												// Trace: src/VX_cache_init.sv:69:5
												wire flush_req_enable = |flush_req_mask;
												// Trace: src/VX_cache_init.sv:70:5
												reg [0:0] lock_released;
												reg [0:0] lock_released_n;
												// Trace: src/VX_cache_init.sv:71:5
												reg [0:0] flush_uuid_r;
												reg [0:0] flush_uuid_n;
												// Trace: src/VX_cache_init.sv:72:5
												genvar _gv_i_216;
												for (_gv_i_216 = 0; _gv_i_216 < NUM_REQS; _gv_i_216 = _gv_i_216 + 1) begin : g_core_bus_out_req
													localparam i = _gv_i_216;
													// Trace: src/VX_cache_init.sv:73:9
													wire input_enable = ~flush_req_enable || lock_released[i];
													// Trace: src/VX_cache_init.sv:74:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_valid && input_enable;
													// Trace: src/VX_cache_init.sv:75:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_data;
													// Trace: src/VX_cache_init.sv:76:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_ready && input_enable;
												end
												// Trace: src/VX_cache_init.sv:78:5
												genvar _gv_i_217;
												for (_gv_i_217 = 0; _gv_i_217 < NUM_REQS; _gv_i_217 = _gv_i_217 + 1) begin : g_core_bus_in_rsp
													localparam i = _gv_i_217;
													// Trace: src/VX_cache_init.sv:79:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].rsp_valid;
													// Trace: src/VX_cache_init.sv:80:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].rsp_data;
													// Trace: src/VX_cache_init.sv:81:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].rsp_ready;
												end
												// Trace: src/VX_cache_init.sv:83:5
												reg [0:0] core_bus_out_uuid;
												// Trace: src/VX_cache_init.sv:84:5
												wire [0:0] core_bus_out_ready;
												// Trace: src/VX_cache_init.sv:85:5
												genvar _gv_i_218;
												for (_gv_i_218 = 0; _gv_i_218 < NUM_REQS; _gv_i_218 = _gv_i_218 + 1) begin : g_core_bus_out_uuid
													localparam i = _gv_i_218;
													if (1) begin : g_uuid
														// Trace: src/VX_cache_init.sv:87:13
														wire [1:1] sv2v_tmp_EFEFC;
														assign sv2v_tmp_EFEFC = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_data[2-:1];
														always @(*) core_bus_out_uuid[i+:1] = sv2v_tmp_EFEFC;
													end
												end
												// Trace: src/VX_cache_init.sv:92:5
												genvar _gv_i_219;
												for (_gv_i_219 = 0; _gv_i_219 < NUM_REQS; _gv_i_219 = _gv_i_219 + 1) begin : g_core_bus_out_ready
													localparam i = _gv_i_219;
													// Trace: src/VX_cache_init.sv:93:9
													assign core_bus_out_ready[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_ready;
												end
												// Trace: src/VX_cache_init.sv:95:5
												always @(*) begin
													// Trace: src/VX_cache_init.sv:96:9
													state_n = state;
													// Trace: src/VX_cache_init.sv:97:9
													flush_done_n = flush_done;
													// Trace: src/VX_cache_init.sv:98:9
													lock_released_n = lock_released;
													// Trace: src/VX_cache_init.sv:99:9
													flush_uuid_n = flush_uuid_r;
													// Trace: src/VX_cache_init.sv:100:9
													case (state)
														default:
															// Trace: src/VX_cache_init.sv:102:17
															if (flush_req_enable) begin
																// Trace: src/VX_cache_init.sv:103:21
																state_n = STATE_FLUSH;
																// Trace: src/VX_cache_init.sv:104:21
																begin : sv2v_autoblock_1
																	// Trace: src/VX_cache_init.sv:104:26
																	integer i;
																	// Trace: src/VX_cache_init.sv:104:26
																	for (i = 0; i >= 0; i = i - 1)
																		begin
																			// Trace: src/VX_cache_init.sv:105:25
																			if (flush_req_mask[i])
																				// Trace: src/VX_cache_init.sv:106:29
																				flush_uuid_n = core_bus_out_uuid[i+:1];
																		end
																end
															end
														STATE_WAIT1:
															// Trace: src/VX_cache_init.sv:112:17
															if (no_inflight_reqs)
																// Trace: src/VX_cache_init.sv:113:21
																state_n = STATE_FLUSH;
														STATE_FLUSH:
															// Trace: src/VX_cache_init.sv:117:17
															state_n = STATE_WAIT2;
														STATE_WAIT2: begin
															// Trace: src/VX_cache_init.sv:120:17
															flush_done_n = flush_done | flush_end;
															// Trace: src/VX_cache_init.sv:121:17
															if (flush_done_n == {NUM_BANKS {1'b1}}) begin
																// Trace: src/VX_cache_init.sv:122:21
																state_n = STATE_DONE;
																// Trace: src/VX_cache_init.sv:123:21
																flush_done_n = 1'sb0;
																// Trace: src/VX_cache_init.sv:124:21
																lock_released_n = flush_req_mask;
															end
														end
														STATE_DONE: begin
															// Trace: src/VX_cache_init.sv:128:17
															lock_released_n = lock_released & ~core_bus_out_ready;
															// Trace: src/VX_cache_init.sv:129:17
															if (lock_released_n == 0)
																// Trace: src/VX_cache_init.sv:130:21
																state_n = STATE_IDLE;
														end
													endcase
												end
												// Trace: src/VX_cache_init.sv:135:5
												always @(posedge clk) begin
													// Trace: src/VX_cache_init.sv:136:9
													if (reset) begin
														// Trace: src/VX_cache_init.sv:137:13
														state <= STATE_IDLE;
														// Trace: src/VX_cache_init.sv:138:13
														flush_done <= 1'sb0;
														// Trace: src/VX_cache_init.sv:139:13
														lock_released <= 1'sb0;
													end
													else begin
														// Trace: src/VX_cache_init.sv:141:13
														state <= state_n;
														// Trace: src/VX_cache_init.sv:142:13
														flush_done <= flush_done_n;
														// Trace: src/VX_cache_init.sv:143:13
														lock_released <= lock_released_n;
													end
													// Trace: src/VX_cache_init.sv:145:9
													flush_uuid_r <= flush_uuid_n;
												end
												// Trace: src/VX_cache_init.sv:147:5
												assign flush_begin = {NUM_BANKS {state == STATE_FLUSH}};
												// Trace: src/VX_cache_init.sv:148:5
												assign flush_uuid = flush_uuid_r;
											end
											assign cache_init.clk = clk;
											assign cache_init.reset = reset;
											assign cache_init.bank_req_fire = per_bank_core_req_fire;
											assign per_bank_flush_begin = cache_init.flush_begin;
											assign flush_uuid = cache_init.flush_uuid;
											assign cache_init.flush_end = per_bank_flush_end;
											// Trace: src/VX_cache.sv:73:5
											// expanded interface instance: mem_bus_tmp_if
											localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
											localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH;
											genvar _arr_4FE36;
											for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [610:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [516:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache.sv:77:5
											wire [0:0] mem_rsp_queue_valid;
											// Trace: src/VX_cache.sv:78:5
											wire [516:0] mem_rsp_queue_data;
											// Trace: src/VX_cache.sv:79:5
											wire [0:0] mem_rsp_queue_ready;
											// Trace: src/VX_cache.sv:80:5
											genvar _gv_i_228;
											for (_gv_i_228 = 0; _gv_i_228 < MEM_PORTS; _gv_i_228 = _gv_i_228 + 1) begin : g_mem_rsp_queue
												localparam i = _gv_i_228;
												// Trace: src/VX_cache.sv:81:9
												VX_elastic_buffer #(
													.DATAW(MEM_RSP_DATAW),
													.SIZE(MRSQ_SIZE),
													.OUT_REG(1'd0)
												) mem_rsp_queue(
													.clk(clk),
													.reset(reset),
													.valid_in(mem_bus_tmp_if[i].rsp_valid),
													.data_in(mem_bus_tmp_if[i].rsp_data),
													.ready_in(mem_bus_tmp_if[i].rsp_ready),
													.valid_out(mem_rsp_queue_valid[i]),
													.data_out(mem_rsp_queue_data[i * 517+:517]),
													.ready_out(mem_rsp_queue_ready[i])
												);
											end
											// Trace: src/VX_cache.sv:96:5
											wire [516:0] mem_rsp_queue_data_s;
											// Trace: src/VX_cache.sv:97:5
											wire [0:0] mem_rsp_queue_sel;
											// Trace: src/VX_cache.sv:98:5
											genvar _gv_i_229;
											for (_gv_i_229 = 0; _gv_i_229 < MEM_PORTS; _gv_i_229 = _gv_i_229 + 1) begin : g_mem_rsp_queue_data_s
												localparam i = _gv_i_229;
												// Trace: src/VX_cache.sv:99:9
												wire [4:0] mem_rsp_tag_s = mem_rsp_queue_data[(i * 517) + 4-:5];
												// Trace: src/VX_cache.sv:100:9
												wire [511:0] mem_rsp_data_s = mem_rsp_queue_data[(i * 517) + 516-:512];
												// Trace: src/VX_cache.sv:101:9
												assign mem_rsp_queue_data_s[i * 517+:517] = {mem_rsp_data_s, mem_rsp_tag_s};
											end
											// Trace: src/VX_cache.sv:103:5
											genvar _gv_i_230;
											for (_gv_i_230 = 0; _gv_i_230 < MEM_PORTS; _gv_i_230 = _gv_i_230 + 1) begin : g_mem_rsp_queue_sel
												localparam i = _gv_i_230;
												if (1) begin : g_singlebank
													// Trace: src/VX_cache.sv:118:13
													assign mem_rsp_queue_sel[i+:1] = 0;
												end
											end
											// Trace: src/VX_cache.sv:121:5
											wire [0:0] per_bank_mem_rsp_valid;
											// Trace: src/VX_cache.sv:122:5
											wire [516:0] per_bank_mem_rsp_pdata;
											// Trace: src/VX_cache.sv:123:5
											wire [0:0] per_bank_mem_rsp_ready;
											// Trace: src/VX_cache.sv:124:5
											VX_stream_omega #(
												.NUM_INPUTS(MEM_PORTS),
												.NUM_OUTPUTS(NUM_BANKS),
												.DATAW(517),
												.ARBITER("R"),
												.OUT_BUF(3)
											) mem_rsp_xbar(
												.clk(clk),
												.reset(reset),
												.valid_in(mem_rsp_queue_valid),
												.data_in(mem_rsp_queue_data_s),
												.sel_in(mem_rsp_queue_sel),
												.ready_in(mem_rsp_queue_ready),
												.valid_out(per_bank_mem_rsp_valid),
												.data_out(per_bank_mem_rsp_pdata),
												.sel_out(),
												.ready_out(per_bank_mem_rsp_ready),
												.collisions()
											);
											// Trace: src/VX_cache.sv:143:5
											wire [511:0] per_bank_mem_rsp_data;
											// Trace: src/VX_cache.sv:144:5
											wire [4:0] per_bank_mem_rsp_tag;
											// Trace: src/VX_cache.sv:145:5
											genvar _gv_i_231;
											for (_gv_i_231 = 0; _gv_i_231 < NUM_BANKS; _gv_i_231 = _gv_i_231 + 1) begin : g_per_bank_mem_rsp_data
												localparam i = _gv_i_231;
												// Trace: src/VX_cache.sv:146:9
												assign {per_bank_mem_rsp_data[i * 512+:512], per_bank_mem_rsp_tag[i * 5+:5]} = per_bank_mem_rsp_pdata[i * 517+:517];
											end
											// Trace: src/VX_cache.sv:151:5
											wire [0:0] per_bank_core_req_valid;
											// Trace: src/VX_cache.sv:152:5
											wire [25:0] per_bank_core_req_addr;
											// Trace: src/VX_cache.sv:153:5
											wire [0:0] per_bank_core_req_rw;
											// Trace: src/VX_cache.sv:154:5
											wire [3:0] per_bank_core_req_wsel;
											// Trace: src/VX_cache.sv:155:5
											wire [3:0] per_bank_core_req_byteen;
											// Trace: src/VX_cache.sv:156:5
											wire [31:0] per_bank_core_req_data;
											// Trace: src/VX_cache.sv:157:5
											wire [2:0] per_bank_core_req_tag;
											// Trace: src/VX_cache.sv:158:5
											wire [0:0] per_bank_core_req_idx;
											// Trace: src/VX_cache.sv:159:5
											wire [2:0] per_bank_core_req_flags;
											// Trace: src/VX_cache.sv:160:5
											wire [0:0] per_bank_core_req_ready;
											// Trace: src/VX_cache.sv:161:5
											wire [0:0] per_bank_core_rsp_valid;
											// Trace: src/VX_cache.sv:162:5
											wire [31:0] per_bank_core_rsp_data;
											// Trace: src/VX_cache.sv:163:5
											wire [2:0] per_bank_core_rsp_tag;
											// Trace: src/VX_cache.sv:164:5
											wire [0:0] per_bank_core_rsp_idx;
											// Trace: src/VX_cache.sv:165:5
											wire [0:0] per_bank_core_rsp_ready;
											// Trace: src/VX_cache.sv:166:5
											wire [0:0] per_bank_mem_req_valid;
											// Trace: src/VX_cache.sv:167:5
											wire [25:0] per_bank_mem_req_addr;
											// Trace: src/VX_cache.sv:168:5
											wire [0:0] per_bank_mem_req_rw;
											// Trace: src/VX_cache.sv:169:5
											wire [63:0] per_bank_mem_req_byteen;
											// Trace: src/VX_cache.sv:170:5
											wire [511:0] per_bank_mem_req_data;
											// Trace: src/VX_cache.sv:171:5
											wire [4:0] per_bank_mem_req_tag;
											// Trace: src/VX_cache.sv:172:5
											wire [2:0] per_bank_mem_req_flags;
											// Trace: src/VX_cache.sv:173:5
											wire [0:0] per_bank_mem_req_ready;
											// Trace: src/VX_cache.sv:174:5
											wire [0:0] core_req_valid;
											// Trace: src/VX_cache.sv:175:5
											wire [29:0] core_req_addr;
											// Trace: src/VX_cache.sv:176:5
											wire [0:0] core_req_rw;
											// Trace: src/VX_cache.sv:177:5
											wire [3:0] core_req_byteen;
											// Trace: src/VX_cache.sv:178:5
											wire [31:0] core_req_data;
											// Trace: src/VX_cache.sv:179:5
											wire [2:0] core_req_tag;
											// Trace: src/VX_cache.sv:180:5
											wire [2:0] core_req_flags;
											// Trace: src/VX_cache.sv:181:5
											wire [0:0] core_req_ready;
											// Trace: src/VX_cache.sv:182:5
											wire [25:0] core_req_line_addr;
											// Trace: src/VX_cache.sv:183:5
											wire [0:0] core_req_bid;
											// Trace: src/VX_cache.sv:184:5
											wire [3:0] core_req_wsel;
											// Trace: src/VX_cache.sv:185:5
											wire [72:0] core_req_data_in;
											// Trace: src/VX_cache.sv:186:5
											wire [72:0] core_req_data_out;
											// Trace: src/VX_cache.sv:187:5
											genvar _gv_i_232;
											for (_gv_i_232 = 0; _gv_i_232 < NUM_REQS; _gv_i_232 = _gv_i_232 + 1) begin : g_core_req
												localparam i = _gv_i_232;
												// Trace: src/VX_cache.sv:188:9
												assign core_req_valid[i] = core_bus2_if[i].req_valid;
												// Trace: src/VX_cache.sv:189:9
												assign core_req_rw[i] = core_bus2_if[i].req_data[72];
												// Trace: src/VX_cache.sv:190:9
												assign core_req_byteen[i * 4+:4] = core_bus2_if[i].req_data[9-:4];
												// Trace: src/VX_cache.sv:191:9
												assign core_req_addr[i * 30+:30] = core_bus2_if[i].req_data[71-:30];
												// Trace: src/VX_cache.sv:192:9
												assign core_req_data[i * 32+:32] = core_bus2_if[i].req_data[41-:32];
												// Trace: src/VX_cache.sv:193:9
												assign core_req_tag[i * 3+:3] = core_bus2_if[i].req_data[2-:3];
												// Trace: src/VX_cache.sv:194:9
												assign core_req_flags[i * 3+:3] = sv2v_cast_3(core_bus2_if[i].req_data[5-:3]);
												// Trace: src/VX_cache.sv:195:9
												assign core_bus2_if[i].req_ready = core_req_ready[i];
											end
											// Trace: src/VX_cache.sv:197:5
											genvar _gv_i_233;
											for (_gv_i_233 = 0; _gv_i_233 < NUM_REQS; _gv_i_233 = _gv_i_233 + 1) begin : g_core_req_wsel
												localparam i = _gv_i_233;
												if (1) begin : g_wsel
													// Trace: src/VX_cache.sv:199:13
													assign core_req_wsel[i * 4+:4] = core_req_addr[i * 30+:WORD_SEL_BITS];
												end
											end
											// Trace: src/VX_cache.sv:204:5
											genvar _gv_i_234;
											for (_gv_i_234 = 0; _gv_i_234 < NUM_REQS; _gv_i_234 = _gv_i_234 + 1) begin : g_core_req_line_addr
												localparam i = _gv_i_234;
												// Trace: src/VX_cache.sv:205:9
												assign core_req_line_addr[i * 26+:26] = core_req_addr[(i * 30) + 4+:LINE_ADDR_WIDTH];
											end
											// Trace: src/VX_cache.sv:207:5
											genvar _gv_i_235;
											for (_gv_i_235 = 0; _gv_i_235 < NUM_REQS; _gv_i_235 = _gv_i_235 + 1) begin : g_core_req_bid
												localparam i = _gv_i_235;
												if (1) begin : g_singlebank
													// Trace: src/VX_cache.sv:211:13
													assign core_req_bid[i+:1] = 1'sb0;
												end
											end
											// Trace: src/VX_cache.sv:214:5
											genvar _gv_i_236;
											for (_gv_i_236 = 0; _gv_i_236 < NUM_REQS; _gv_i_236 = _gv_i_236 + 1) begin : g_core_req_data_in
												localparam i = _gv_i_236;
												// Trace: src/VX_cache.sv:215:9
												assign core_req_data_in[i * 73+:73] = {core_req_line_addr[i * 26+:26], core_req_rw[i], core_req_wsel[i * 4+:4], core_req_byteen[i * 4+:4], core_req_data[i * 32+:32], core_req_tag[i * 3+:3], core_req_flags[i * 3+:3]};
											end
											// Trace: src/VX_cache.sv:225:5
											assign per_bank_core_req_fire = per_bank_core_req_valid & per_bank_mem_req_ready;
											// Trace: src/VX_cache.sv:226:5
											localparam VX_gpu_pkg_PERF_CTR_BITS = 44;
											VX_stream_xbar #(
												.NUM_INPUTS(NUM_REQS),
												.NUM_OUTPUTS(NUM_BANKS),
												.DATAW(CORE_REQ_DATAW),
												.PERF_CTR_BITS(VX_gpu_pkg_PERF_CTR_BITS),
												.ARBITER("R"),
												.OUT_BUF(REQ_XBAR_BUF)
											) core_req_xbar(
												.clk(clk),
												.reset(reset),
												.collisions(),
												.valid_in(core_req_valid),
												.data_in(core_req_data_in),
												.sel_in(core_req_bid),
												.ready_in(core_req_ready),
												.valid_out(per_bank_core_req_valid),
												.data_out(core_req_data_out),
												.sel_out(per_bank_core_req_idx),
												.ready_out(per_bank_core_req_ready)
											);
											// Trace: src/VX_cache.sv:246:5
											genvar _gv_i_237;
											for (_gv_i_237 = 0; _gv_i_237 < NUM_BANKS; _gv_i_237 = _gv_i_237 + 1) begin : g_core_req_data_out
												localparam i = _gv_i_237;
												// Trace: src/VX_cache.sv:247:9
												assign {per_bank_core_req_addr[i * 26+:26], per_bank_core_req_rw[i], per_bank_core_req_wsel[i * 4+:4], per_bank_core_req_byteen[i * 4+:4], per_bank_core_req_data[i * 32+:32], per_bank_core_req_tag[i * 3+:3], per_bank_core_req_flags[i * 3+:3]} = core_req_data_out[i * 73+:73];
											end
											// Trace: src/VX_cache.sv:257:5
											genvar _gv_bank_id_1;
											for (_gv_bank_id_1 = 0; _gv_bank_id_1 < NUM_BANKS; _gv_bank_id_1 = _gv_bank_id_1 + 1) begin : g_banks
												localparam bank_id = _gv_bank_id_1;
												// Trace: src/VX_cache.sv:258:9
												VX_cache_bank #(
													.BANK_ID(bank_id),
													.INSTANCE_ID(""),
													.CACHE_SIZE(CACHE_SIZE),
													.LINE_SIZE(LINE_SIZE),
													.NUM_BANKS(NUM_BANKS),
													.NUM_WAYS(NUM_WAYS),
													.WORD_SIZE(WORD_SIZE),
													.NUM_REQS(NUM_REQS),
													.WRITE_ENABLE(WRITE_ENABLE),
													.WRITEBACK(WRITEBACK),
													.DIRTY_BYTES(DIRTY_BYTES),
													.REPL_POLICY(REPL_POLICY),
													.CRSQ_SIZE(CRSQ_SIZE),
													.MSHR_SIZE(MSHR_SIZE),
													.MREQ_SIZE(MREQ_SIZE),
													.TAG_WIDTH(TAG_WIDTH),
													.CORE_OUT_REG((CORE_RSP_BUF_ENABLE ? 0 : ((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : (CORE_OUT_BUF & 7) - 2))),
													.MEM_OUT_REG((MEM_REQ_BUF_ENABLE ? 0 : ((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : (MEM_OUT_BUF & 7) - 2)))
												) bank(
													.clk(clk),
													.reset(reset),
													.core_req_valid(per_bank_core_req_valid[bank_id]),
													.core_req_addr(per_bank_core_req_addr[bank_id * 26+:26]),
													.core_req_rw(per_bank_core_req_rw[bank_id]),
													.core_req_wsel(per_bank_core_req_wsel[bank_id * 4+:4]),
													.core_req_byteen(per_bank_core_req_byteen[bank_id * 4+:4]),
													.core_req_data(per_bank_core_req_data[bank_id * 32+:32]),
													.core_req_tag(per_bank_core_req_tag[bank_id * 3+:3]),
													.core_req_idx(per_bank_core_req_idx[bank_id+:1]),
													.core_req_flags(per_bank_core_req_flags[bank_id * 3+:3]),
													.core_req_ready(per_bank_core_req_ready[bank_id]),
													.core_rsp_valid(per_bank_core_rsp_valid[bank_id]),
													.core_rsp_data(per_bank_core_rsp_data[bank_id * 32+:32]),
													.core_rsp_tag(per_bank_core_rsp_tag[bank_id * 3+:3]),
													.core_rsp_idx(per_bank_core_rsp_idx[bank_id+:1]),
													.core_rsp_ready(per_bank_core_rsp_ready[bank_id]),
													.mem_req_valid(per_bank_mem_req_valid[bank_id]),
													.mem_req_addr(per_bank_mem_req_addr[bank_id * 26+:26]),
													.mem_req_rw(per_bank_mem_req_rw[bank_id]),
													.mem_req_byteen(per_bank_mem_req_byteen[bank_id * 64+:64]),
													.mem_req_data(per_bank_mem_req_data[bank_id * 512+:512]),
													.mem_req_tag(per_bank_mem_req_tag[bank_id * 5+:5]),
													.mem_req_flags(per_bank_mem_req_flags[bank_id * 3+:3]),
													.mem_req_ready(per_bank_mem_req_ready[bank_id]),
													.mem_rsp_valid(per_bank_mem_rsp_valid[bank_id]),
													.mem_rsp_data(per_bank_mem_rsp_data[bank_id * 512+:512]),
													.mem_rsp_tag(per_bank_mem_rsp_tag[bank_id * 5+:5]),
													.mem_rsp_ready(per_bank_mem_rsp_ready[bank_id]),
													.flush_begin(per_bank_flush_begin[bank_id]),
													.flush_uuid(flush_uuid),
													.flush_end(per_bank_flush_end[bank_id])
												);
											end
											// Trace: src/VX_cache.sv:312:5
											wire [34:0] core_rsp_data_in;
											// Trace: src/VX_cache.sv:313:5
											wire [34:0] core_rsp_data_out;
											// Trace: src/VX_cache.sv:314:5
											wire [0:0] core_rsp_valid_s;
											// Trace: src/VX_cache.sv:315:5
											wire [31:0] core_rsp_data_s;
											// Trace: src/VX_cache.sv:316:5
											wire [2:0] core_rsp_tag_s;
											// Trace: src/VX_cache.sv:317:5
											wire [0:0] core_rsp_ready_s;
											// Trace: src/VX_cache.sv:318:5
											genvar _gv_i_238;
											for (_gv_i_238 = 0; _gv_i_238 < NUM_BANKS; _gv_i_238 = _gv_i_238 + 1) begin : g_core_rsp_data_in
												localparam i = _gv_i_238;
												// Trace: src/VX_cache.sv:319:9
												assign core_rsp_data_in[i * 35+:35] = {per_bank_core_rsp_data[i * 32+:32], per_bank_core_rsp_tag[i * 3+:3]};
											end
											// Trace: src/VX_cache.sv:321:5
											VX_stream_xbar #(
												.NUM_INPUTS(NUM_BANKS),
												.NUM_OUTPUTS(NUM_REQS),
												.DATAW(CORE_RSP_DATAW),
												.ARBITER("R")
											) core_rsp_xbar(
												.clk(clk),
												.reset(reset),
												.collisions(),
												.valid_in(per_bank_core_rsp_valid),
												.data_in(core_rsp_data_in),
												.sel_in(per_bank_core_rsp_idx),
												.ready_in(per_bank_core_rsp_ready),
												.valid_out(core_rsp_valid_s),
												.data_out(core_rsp_data_out),
												.ready_out(core_rsp_ready_s),
												.sel_out()
											);
											// Trace: src/VX_cache.sv:339:5
											genvar _gv_i_239;
											for (_gv_i_239 = 0; _gv_i_239 < NUM_REQS; _gv_i_239 = _gv_i_239 + 1) begin : g_core_rsp_data_s
												localparam i = _gv_i_239;
												// Trace: src/VX_cache.sv:340:9
												assign {core_rsp_data_s[i * 32+:32], core_rsp_tag_s[i * 3+:3]} = core_rsp_data_out[i * 35+:35];
											end
											// Trace: src/VX_cache.sv:342:5
											genvar _gv_i_240;
											for (_gv_i_240 = 0; _gv_i_240 < NUM_REQS; _gv_i_240 = _gv_i_240 + 1) begin : g_core_rsp_buf
												localparam i = _gv_i_240;
												// Trace: src/VX_cache.sv:343:9
												VX_elastic_buffer #(
													.DATAW(35),
													.SIZE((CORE_RSP_BUF_ENABLE ? ((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : 2) : 0)),
													.OUT_REG(((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : (CORE_OUT_BUF & 7) - 2))
												) core_rsp_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(core_rsp_valid_s[i]),
													.ready_in(core_rsp_ready_s[i]),
													.data_in({core_rsp_data_s[i * 32+:32], core_rsp_tag_s[i * 3+:3]}),
													.data_out({core_bus2_if[i].rsp_data[34-:32], core_bus2_if[i].rsp_data[2-:3]}),
													.valid_out(core_bus2_if[i].rsp_valid),
													.ready_out(core_bus2_if[i].rsp_ready)
												);
											end
											// Trace: src/VX_cache.sv:358:5
											wire [610:0] per_bank_mem_req_pdata;
											// Trace: src/VX_cache.sv:359:5
											genvar _gv_i_241;
											for (_gv_i_241 = 0; _gv_i_241 < NUM_BANKS; _gv_i_241 = _gv_i_241 + 1) begin : g_per_bank_mem_req_pdata
												localparam i = _gv_i_241;
												// Trace: src/VX_cache.sv:360:9
												assign per_bank_mem_req_pdata[i * 611+:611] = {per_bank_mem_req_rw[i], per_bank_mem_req_addr[i * 26+:26], per_bank_mem_req_data[i * 512+:512], per_bank_mem_req_byteen[i * 64+:64], per_bank_mem_req_flags[i * 3+:3], per_bank_mem_req_tag[i * 5+:5]};
											end
											// Trace: src/VX_cache.sv:369:5
											wire [0:0] mem_req_valid;
											// Trace: src/VX_cache.sv:370:5
											wire [610:0] mem_req_pdata;
											// Trace: src/VX_cache.sv:371:5
											wire [0:0] mem_req_ready;
											// Trace: src/VX_cache.sv:372:5
											wire [0:0] mem_req_sel_out;
											// Trace: src/VX_cache.sv:373:5
											VX_stream_arb #(
												.NUM_INPUTS(NUM_BANKS),
												.NUM_OUTPUTS(MEM_PORTS),
												.DATAW(MEM_REQ_DATAW),
												.ARBITER("R")
											) mem_req_arb(
												.clk(clk),
												.reset(reset),
												.valid_in(per_bank_mem_req_valid),
												.data_in(per_bank_mem_req_pdata),
												.ready_in(per_bank_mem_req_ready),
												.valid_out(mem_req_valid),
												.data_out(mem_req_pdata),
												.ready_out(mem_req_ready),
												.sel_out(mem_req_sel_out)
											);
											// Trace: src/VX_cache.sv:389:5
											genvar _gv_i_242;
											for (_gv_i_242 = 0; _gv_i_242 < MEM_PORTS; _gv_i_242 = _gv_i_242 + 1) begin : g_mem_req_buf
												localparam i = _gv_i_242;
												// Trace: src/VX_cache.sv:390:9
												wire mem_req_rw;
												// Trace: src/VX_cache.sv:391:9
												wire [25:0] mem_req_addr;
												// Trace: src/VX_cache.sv:392:9
												wire [511:0] mem_req_data;
												// Trace: src/VX_cache.sv:393:9
												wire [63:0] mem_req_byteen;
												// Trace: src/VX_cache.sv:394:9
												wire [2:0] mem_req_flags;
												// Trace: src/VX_cache.sv:395:9
												wire [4:0] mem_req_tag;
												// Trace: src/VX_cache.sv:396:9
												assign {mem_req_rw, mem_req_addr, mem_req_data, mem_req_byteen, mem_req_flags, mem_req_tag} = mem_req_pdata[i * 611+:611];
												// Trace: src/VX_cache.sv:404:9
												wire [25:0] mem_req_addr_w;
												// Trace: src/VX_cache.sv:405:9
												wire [4:0] mem_req_tag_w;
												// Trace: src/VX_cache.sv:406:9
												wire [2:0] mem_req_flags_w;
												if (1) begin : g_mem_req_tag
													// Trace: src/VX_cache.sv:425:13
													assign mem_req_addr_w = mem_req_addr;
													// Trace: src/VX_cache.sv:426:13
													assign mem_req_tag_w = mem_req_tag;
												end
												// Trace: src/VX_cache.sv:428:9
												VX_elastic_buffer #(
													.DATAW(611),
													.SIZE((MEM_REQ_BUF_ENABLE ? ((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : 2) : 0)),
													.OUT_REG(((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : (MEM_OUT_BUF & 7) - 2))
												) mem_req_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(mem_req_valid[i]),
													.ready_in(mem_req_ready[i]),
													.data_in({mem_req_rw, mem_req_byteen, mem_req_addr_w, mem_req_data, mem_req_tag_w, mem_req_flags}),
													.data_out({mem_bus_tmp_if[i].req_data[610], mem_bus_tmp_if[i].req_data[71-:64], mem_bus_tmp_if[i].req_data[609-:26], mem_bus_tmp_if[i].req_data[583-:512], mem_bus_tmp_if[i].req_data[4-:5], mem_req_flags_w}),
													.valid_out(mem_bus_tmp_if[i].req_valid),
													.ready_out(mem_bus_tmp_if[i].req_ready)
												);
												if (1) begin : g_mem_req_flags
													// Trace: src/VX_cache.sv:443:13
													assign mem_bus_tmp_if[i].req_data[7-:3] = mem_req_flags_w;
												end
												if (WRITE_ENABLE) begin : g_mem_bus_if
													// Trace: src/VX_cache.sv:448:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
													// Trace: src/VX_cache.sv:449:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[i].req_data;
													// Trace: src/VX_cache.sv:450:5
													assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_ready;
													// Trace: src/VX_cache.sv:451:5
													assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_valid;
													// Trace: src/VX_cache.sv:452:5
													assign mem_bus_tmp_if[i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_data;
													// Trace: src/VX_cache.sv:453:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
												end
												else begin : g_mem_bus_if_ro
													// Trace: src/VX_cache.sv:455:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
													// Trace: src/VX_cache.sv:456:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[610] = 0;
													// Trace: src/VX_cache.sv:457:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[609-:26] = mem_bus_tmp_if[i].req_data[609-:26];
													// Trace: src/VX_cache.sv:458:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[583-:512] = 1'sb0;
													// Trace: src/VX_cache.sv:459:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[71-:64] = 1'sb1;
													// Trace: src/VX_cache.sv:460:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[7-:3] = mem_bus_tmp_if[i].req_data[7-:3];
													// Trace: src/VX_cache.sv:461:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[4-:5] = mem_bus_tmp_if[i].req_data[4-:5];
													// Trace: src/VX_cache.sv:462:5
													assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_ready;
													// Trace: src/VX_cache.sv:463:5
													assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_valid;
													// Trace: src/VX_cache.sv:464:5
													assign mem_bus_tmp_if[i].rsp_data[516-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_data[516-:512];
													// Trace: src/VX_cache.sv:465:5
													assign mem_bus_tmp_if[i].rsp_data[4-:5] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_data[4-:5];
													// Trace: src/VX_cache.sv:466:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
												end
											end
										end
										assign cache.clk = clk;
										assign cache.reset = reset;
									end
								end
								assign cache_wrap.clk = clk;
								assign cache_wrap.reset = reset;
							end
							// Trace: src/VX_cache_cluster.sv:120:5
							genvar _gv_i_193;
							for (_gv_i_193 = 0; _gv_i_193 < MEM_PORTS; _gv_i_193 = _gv_i_193 + 1) begin : g_mem_bus_if
								localparam i = _gv_i_193;
								// Trace: src/VX_cache_cluster.sv:121:9
								// expanded interface instance: arb_core_bus_tmp_if
								localparam _param_E788B_DATA_SIZE = LINE_SIZE;
								localparam _param_E788B_TAG_WIDTH = MEM_TAG_WIDTH;
								genvar _arr_E788B;
								for (_arr_E788B = 0; _arr_E788B <= 0; _arr_E788B = _arr_E788B + 1) begin : arb_core_bus_tmp_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_E788B_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_E788B_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:8:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:12:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:20:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:24:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire [610:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire [516:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:30:5
									// Trace: src/VX_mem_bus_if.sv:38:5
								end
								// Trace: src/VX_cache_cluster.sv:125:9
								// expanded interface instance: mem_bus_tmp_if
								localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
								localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH + 0;
								genvar _arr_4FE36;
								for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:8:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:12:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:20:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:24:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire [610:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire [516:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:30:5
									// Trace: src/VX_mem_bus_if.sv:38:5
								end
								genvar _gv_j_20;
								for (_gv_j_20 = 0; _gv_j_20 < NUM_CACHES; _gv_j_20 = _gv_j_20 + 1) begin : g_arb_core_bus_tmp_if
									localparam j = _gv_j_20;
									// Trace: src/VX_cache_cluster.sv:130:5
									assign arb_core_bus_tmp_if[j].req_valid = cache_mem_bus_if[(j * MEM_PORTS) + i].req_valid;
									// Trace: src/VX_cache_cluster.sv:131:5
									assign arb_core_bus_tmp_if[j].req_data = cache_mem_bus_if[(j * MEM_PORTS) + i].req_data;
									// Trace: src/VX_cache_cluster.sv:132:5
									assign cache_mem_bus_if[(j * MEM_PORTS) + i].req_ready = arb_core_bus_tmp_if[j].req_ready;
									// Trace: src/VX_cache_cluster.sv:133:5
									assign cache_mem_bus_if[(j * MEM_PORTS) + i].rsp_valid = arb_core_bus_tmp_if[j].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:134:5
									assign cache_mem_bus_if[(j * MEM_PORTS) + i].rsp_data = arb_core_bus_tmp_if[j].rsp_data;
									// Trace: src/VX_cache_cluster.sv:135:5
									assign arb_core_bus_tmp_if[j].rsp_ready = cache_mem_bus_if[(j * MEM_PORTS) + i].rsp_ready;
								end
								// Trace: src/VX_cache_cluster.sv:137:9
								// expanded module instance: mem_arb
								localparam _bbase_7277A_bus_in_if = 0;
								localparam _bbase_7277A_bus_out_if = 0;
								localparam _param_7277A_NUM_INPUTS = NUM_CACHES;
								localparam _param_7277A_NUM_OUTPUTS = 1;
								localparam _param_7277A_DATA_SIZE = LINE_SIZE;
								localparam _param_7277A_TAG_WIDTH = MEM_TAG_WIDTH;
								localparam _param_7277A_TAG_SEL_IDX = TAG_SEL_IDX;
								localparam _param_7277A_ARBITER = "R";
								localparam _param_7277A_REQ_OUT_BUF = 0;
								localparam _param_7277A_RSP_OUT_BUF = 0;
								if (1) begin : mem_arb
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_arb.sv:2:15
									localparam NUM_INPUTS = _param_7277A_NUM_INPUTS;
									// Trace: src/VX_mem_arb.sv:3:15
									localparam NUM_OUTPUTS = _param_7277A_NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:4:15
									localparam DATA_SIZE = _param_7277A_DATA_SIZE;
									// Trace: src/VX_mem_arb.sv:5:15
									localparam TAG_WIDTH = _param_7277A_TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:6:15
									localparam TAG_SEL_IDX = _param_7277A_TAG_SEL_IDX;
									// Trace: src/VX_mem_arb.sv:7:15
									localparam REQ_OUT_BUF = _param_7277A_REQ_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:8:15
									localparam RSP_OUT_BUF = _param_7277A_RSP_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:9:15
									localparam ARBITER = _param_7277A_ARBITER;
									// Trace: src/VX_mem_arb.sv:10:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_arb.sv:11:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_arb.sv:12:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_arb.sv:14:5
									wire clk;
									// Trace: src/VX_mem_arb.sv:15:5
									wire reset;
									// Trace: src/VX_mem_arb.sv:16:5
									localparam _mbase_bus_in_if = 0;
									// Trace: src/VX_mem_arb.sv:17:5
									localparam _mbase_bus_out_if = 0;
									// Trace: src/VX_mem_arb.sv:19:5
									localparam DATA_WIDTH = 512;
									// Trace: src/VX_mem_arb.sv:20:5
									localparam LOG_NUM_REQS = 0;
									// Trace: src/VX_mem_arb.sv:21:5
									localparam REQ_DATAW = 606 + TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:22:5
									localparam RSP_DATAW = DATA_WIDTH + TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:23:5
									localparam SEL_COUNT = NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:24:5
									wire [0:0] req_valid_in;
									// Trace: src/VX_mem_arb.sv:25:5
									wire [REQ_DATAW - 1:0] req_data_in;
									// Trace: src/VX_mem_arb.sv:26:5
									wire [0:0] req_ready_in;
									// Trace: src/VX_mem_arb.sv:27:5
									wire [0:0] req_valid_out;
									// Trace: src/VX_mem_arb.sv:28:5
									wire [REQ_DATAW - 1:0] req_data_out;
									// Trace: src/VX_mem_arb.sv:29:5
									wire [0:0] req_sel_out;
									// Trace: src/VX_mem_arb.sv:30:5
									wire [0:0] req_ready_out;
									// Trace: src/VX_mem_arb.sv:31:5
									genvar _gv_i_183;
									for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
										localparam i = _gv_i_183;
										// Trace: src/VX_mem_arb.sv:32:9
										assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].arb_core_bus_tmp_if[i + _mbase_bus_in_if].req_valid;
										// Trace: src/VX_mem_arb.sv:33:9
										assign req_data_in[i * 611+:611] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].arb_core_bus_tmp_if[i + _mbase_bus_in_if].req_data;
										// Trace: src/VX_mem_arb.sv:34:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].arb_core_bus_tmp_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:36:5
									VX_stream_arb #(
										.NUM_INPUTS(NUM_INPUTS),
										.NUM_OUTPUTS(NUM_OUTPUTS),
										.DATAW(REQ_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(REQ_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(req_valid_in),
										.ready_in(req_ready_in),
										.data_in(req_data_in),
										.data_out(req_data_out),
										.sel_out(req_sel_out),
										.valid_out(req_valid_out),
										.ready_out(req_ready_out)
									);
									// Trace: src/VX_mem_arb.sv:53:5
									genvar _gv_i_184;
									for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
										localparam i = _gv_i_184;
										// Trace: src/VX_mem_arb.sv:54:9
										wire [TAG_WIDTH - 1:0] req_tag_out;
										// Trace: src/VX_mem_arb.sv:55:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
										// Trace: src/VX_mem_arb.sv:56:9
										assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[610], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[609-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[583-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[71-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[7-:3], req_tag_out} = req_data_out[i * 611+:611];
										// Trace: src/VX_mem_arb.sv:64:9
										assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
										if (1) begin : g_req_tag_out
											// Trace: src/VX_mem_arb.sv:76:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[4-:5] = req_tag_out;
										end
									end
									// Trace: src/VX_mem_arb.sv:79:5
									wire [0:0] rsp_valid_out;
									// Trace: src/VX_mem_arb.sv:80:5
									wire [RSP_DATAW - 1:0] rsp_data_out;
									// Trace: src/VX_mem_arb.sv:81:5
									wire [0:0] rsp_ready_out;
									// Trace: src/VX_mem_arb.sv:82:5
									wire [0:0] rsp_valid_in;
									// Trace: src/VX_mem_arb.sv:83:5
									wire [RSP_DATAW - 1:0] rsp_data_in;
									// Trace: src/VX_mem_arb.sv:84:5
									wire [0:0] rsp_ready_in;
									// Trace: src/VX_mem_arb.sv:85:5
									if (1) begin : g_rsp_arb
										genvar _gv_i_186;
										for (_gv_i_186 = 0; _gv_i_186 < NUM_OUTPUTS; _gv_i_186 = _gv_i_186 + 1) begin : g_rsp_data_in
											localparam i = _gv_i_186;
											// Trace: src/VX_mem_arb.sv:120:13
											assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
											// Trace: src/VX_mem_arb.sv:121:13
											assign rsp_data_in[i * 517+:517] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
											// Trace: src/VX_mem_arb.sv:122:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
										end
										// Trace: src/VX_mem_arb.sv:124:9
										VX_stream_arb #(
											.NUM_INPUTS(NUM_OUTPUTS),
											.NUM_OUTPUTS(NUM_INPUTS),
											.DATAW(RSP_DATAW),
											.ARBITER(ARBITER),
											.OUT_BUF(RSP_OUT_BUF)
										) req_arb(
											.clk(clk),
											.reset(reset),
											.valid_in(rsp_valid_in),
											.ready_in(rsp_ready_in),
											.data_in(rsp_data_in),
											.data_out(rsp_data_out),
											.valid_out(rsp_valid_out),
											.ready_out(rsp_ready_out),
											.sel_out()
										);
									end
									// Trace: src/VX_mem_arb.sv:142:5
									genvar _gv_i_187;
									for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
										localparam i = _gv_i_187;
										// Trace: src/VX_mem_arb.sv:143:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].arb_core_bus_tmp_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
										// Trace: src/VX_mem_arb.sv:144:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].arb_core_bus_tmp_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 517+:517];
										// Trace: src/VX_mem_arb.sv:145:9
										assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache.g_mem_bus_if[_gv_i_193].arb_core_bus_tmp_if[i + _mbase_bus_in_if].rsp_ready;
									end
								end
								assign mem_arb.clk = clk;
								assign mem_arb.reset = reset;
								if (WRITE_ENABLE) begin : g_we
									// Trace: src/VX_cache_cluster.sv:153:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[0].req_valid;
									// Trace: src/VX_cache_cluster.sv:154:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[0].req_data;
									// Trace: src/VX_cache_cluster.sv:155:5
									assign mem_bus_tmp_if[0].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
									// Trace: src/VX_cache_cluster.sv:156:5
									assign mem_bus_tmp_if[0].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:157:5
									assign mem_bus_tmp_if[0].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
									// Trace: src/VX_cache_cluster.sv:158:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[0].rsp_ready;
								end
								else begin : g_ro
									// Trace: src/VX_cache_cluster.sv:160:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[0].req_valid;
									// Trace: src/VX_cache_cluster.sv:161:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data[610] = 0;
									// Trace: src/VX_cache_cluster.sv:162:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data[609-:26] = mem_bus_tmp_if[0].req_data[609-:26];
									// Trace: src/VX_cache_cluster.sv:163:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data[583-:512] = 1'sb0;
									// Trace: src/VX_cache_cluster.sv:164:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data[71-:64] = 1'sb1;
									// Trace: src/VX_cache_cluster.sv:165:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data[7-:3] = mem_bus_tmp_if[0].req_data[7-:3];
									// Trace: src/VX_cache_cluster.sv:166:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_data[4-:5] = mem_bus_tmp_if[0].req_data[4-:5];
									// Trace: src/VX_cache_cluster.sv:167:5
									assign mem_bus_tmp_if[0].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
									// Trace: src/VX_cache_cluster.sv:168:5
									assign mem_bus_tmp_if[0].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:169:5
									assign mem_bus_tmp_if[0].rsp_data[516-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[516-:512];
									// Trace: src/VX_cache_cluster.sv:170:5
									assign mem_bus_tmp_if[0].rsp_data[4-:5] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[4-:5];
									// Trace: src/VX_cache_cluster.sv:171:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.icache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[0].rsp_ready;
								end
							end
						end
						assign icache.clk = clk;
						assign icache.reset = icache_reset;
						// Trace: src/VX_socket.sv:53:5
						localparam VX_gpu_pkg_DCACHE_MERGED_REQS = 1;
						localparam VX_gpu_pkg_DCACHE_MEM_BATCHES = 1;
						localparam VX_gpu_pkg_DCACHE_TAG_ID_BITS = 2;
						localparam VX_gpu_pkg_DCACHE_TAG_WIDTH = 3;
						// expanded interface instance: per_core_dcache_bus_if
						localparam _param_F6DD5_DATA_SIZE = VX_gpu_pkg_DCACHE_WORD_SIZE;
						localparam _param_F6DD5_TAG_WIDTH = VX_gpu_pkg_DCACHE_TAG_WIDTH;
						genvar _arr_F6DD5;
						for (_arr_F6DD5 = 0; _arr_F6DD5 <= 0; _arr_F6DD5 = _arr_F6DD5 + 1) begin : per_core_dcache_bus_if
							// removed import VX_gpu_pkg::*;
							// Trace: src/VX_mem_bus_if.sv:2:15
							localparam DATA_SIZE = _param_F6DD5_DATA_SIZE;
							// Trace: src/VX_mem_bus_if.sv:3:15
							localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
							localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
							localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
							// Trace: src/VX_mem_bus_if.sv:4:15
							localparam TAG_WIDTH = _param_F6DD5_TAG_WIDTH;
							// Trace: src/VX_mem_bus_if.sv:5:15
							localparam MEM_ADDR_WIDTH = 32;
							// Trace: src/VX_mem_bus_if.sv:6:15
							localparam ADDR_WIDTH = 28;
							// Trace: src/VX_mem_bus_if.sv:8:5
							localparam VX_gpu_pkg_UUID_WIDTH = 1;
							// removed localparam type tag_t
							// Trace: src/VX_mem_bus_if.sv:12:5
							// removed localparam type req_data_t
							// Trace: src/VX_mem_bus_if.sv:20:5
							// removed localparam type rsp_data_t
							// Trace: src/VX_mem_bus_if.sv:24:5
							wire req_valid;
							// Trace: src/VX_mem_bus_if.sv:25:5
							wire [178:0] req_data;
							// Trace: src/VX_mem_bus_if.sv:26:5
							wire req_ready;
							// Trace: src/VX_mem_bus_if.sv:27:5
							wire rsp_valid;
							// Trace: src/VX_mem_bus_if.sv:28:5
							wire [130:0] rsp_data;
							// Trace: src/VX_mem_bus_if.sv:29:5
							wire rsp_ready;
							// Trace: src/VX_mem_bus_if.sv:30:5
							// Trace: src/VX_mem_bus_if.sv:38:5
						end
						// Trace: src/VX_socket.sv:57:5
						localparam VX_gpu_pkg_DCACHE_LINE_SIZE = 64;
						localparam VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH = 6;
						// expanded interface instance: dcache_mem_bus_if
						localparam _param_28DB2_DATA_SIZE = VX_gpu_pkg_DCACHE_LINE_SIZE;
						localparam _param_28DB2_TAG_WIDTH = VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH;
						genvar _arr_28DB2;
						for (_arr_28DB2 = 0; _arr_28DB2 <= 0; _arr_28DB2 = _arr_28DB2 + 1) begin : dcache_mem_bus_if
							// removed import VX_gpu_pkg::*;
							// Trace: src/VX_mem_bus_if.sv:2:15
							localparam DATA_SIZE = _param_28DB2_DATA_SIZE;
							// Trace: src/VX_mem_bus_if.sv:3:15
							localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
							localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
							localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
							// Trace: src/VX_mem_bus_if.sv:4:15
							localparam TAG_WIDTH = _param_28DB2_TAG_WIDTH;
							// Trace: src/VX_mem_bus_if.sv:5:15
							localparam MEM_ADDR_WIDTH = 32;
							// Trace: src/VX_mem_bus_if.sv:6:15
							localparam ADDR_WIDTH = 26;
							// Trace: src/VX_mem_bus_if.sv:8:5
							localparam VX_gpu_pkg_UUID_WIDTH = 1;
							// removed localparam type tag_t
							// Trace: src/VX_mem_bus_if.sv:12:5
							// removed localparam type req_data_t
							// Trace: src/VX_mem_bus_if.sv:20:5
							// removed localparam type rsp_data_t
							// Trace: src/VX_mem_bus_if.sv:24:5
							wire req_valid;
							// Trace: src/VX_mem_bus_if.sv:25:5
							wire [611:0] req_data;
							// Trace: src/VX_mem_bus_if.sv:26:5
							wire req_ready;
							// Trace: src/VX_mem_bus_if.sv:27:5
							wire rsp_valid;
							// Trace: src/VX_mem_bus_if.sv:28:5
							wire [517:0] rsp_data;
							// Trace: src/VX_mem_bus_if.sv:29:5
							wire rsp_ready;
							// Trace: src/VX_mem_bus_if.sv:30:5
							// Trace: src/VX_mem_bus_if.sv:38:5
						end
						// Trace: src/VX_socket.sv:61:5
						wire [0:0] dcache_reset;
						// Trace: src/VX_socket.sv:62:5
						VX_reset_relay #(
							.N(1),
							.MAX_FANOUT(0)
						) __dcache_reset(
							.clk(clk),
							.reset(reset),
							.reset_o(dcache_reset)
						);
						// Trace: src/VX_socket.sv:67:5
						// expanded module instance: dcache
						localparam _bbase_CC492_core_bus_if = 0;
						localparam _bbase_CC492_mem_bus_if = 0;
						localparam _param_CC492_INSTANCE_ID = "";
						localparam _param_CC492_NUM_UNITS = 1;
						localparam _param_CC492_NUM_INPUTS = 1;
						localparam _param_CC492_TAG_SEL_IDX = 0;
						localparam _param_CC492_CACHE_SIZE = 16384;
						localparam _param_CC492_LINE_SIZE = VX_gpu_pkg_DCACHE_LINE_SIZE;
						localparam _param_CC492_NUM_BANKS = VX_gpu_pkg_DCACHE_NUM_REQS;
						localparam _param_CC492_NUM_WAYS = 4;
						localparam _param_CC492_WORD_SIZE = VX_gpu_pkg_DCACHE_WORD_SIZE;
						localparam _param_CC492_NUM_REQS = VX_gpu_pkg_DCACHE_NUM_REQS;
						localparam _param_CC492_MEM_PORTS = VX_gpu_pkg_DCACHE_NUM_REQS;
						localparam _param_CC492_CRSQ_SIZE = 2;
						localparam _param_CC492_MSHR_SIZE = 16;
						localparam _param_CC492_MRSQ_SIZE = 4;
						localparam _param_CC492_MREQ_SIZE = 4;
						localparam _param_CC492_TAG_WIDTH = VX_gpu_pkg_DCACHE_TAG_WIDTH;
						localparam _param_CC492_WRITE_ENABLE = 1;
						localparam _param_CC492_WRITEBACK = 0;
						localparam _param_CC492_DIRTY_BYTES = 0;
						localparam _param_CC492_REPL_POLICY = 1;
						localparam _param_CC492_NC_ENABLE = 1;
						localparam _param_CC492_CORE_OUT_BUF = 3;
						localparam _param_CC492_MEM_OUT_BUF = 2;
						if (1) begin : dcache
							// removed import VX_gpu_pkg::*;
							// Trace: src/VX_cache_cluster.sv:2:15
							localparam INSTANCE_ID = _param_CC492_INSTANCE_ID;
							// Trace: src/VX_cache_cluster.sv:3:15
							localparam NUM_UNITS = _param_CC492_NUM_UNITS;
							// Trace: src/VX_cache_cluster.sv:4:15
							localparam NUM_INPUTS = _param_CC492_NUM_INPUTS;
							// Trace: src/VX_cache_cluster.sv:5:15
							localparam TAG_SEL_IDX = _param_CC492_TAG_SEL_IDX;
							// Trace: src/VX_cache_cluster.sv:6:15
							localparam NUM_REQS = _param_CC492_NUM_REQS;
							// Trace: src/VX_cache_cluster.sv:7:15
							localparam MEM_PORTS = _param_CC492_MEM_PORTS;
							// Trace: src/VX_cache_cluster.sv:8:15
							localparam CACHE_SIZE = _param_CC492_CACHE_SIZE;
							// Trace: src/VX_cache_cluster.sv:9:15
							localparam LINE_SIZE = _param_CC492_LINE_SIZE;
							// Trace: src/VX_cache_cluster.sv:10:15
							localparam NUM_BANKS = _param_CC492_NUM_BANKS;
							// Trace: src/VX_cache_cluster.sv:11:15
							localparam NUM_WAYS = _param_CC492_NUM_WAYS;
							// Trace: src/VX_cache_cluster.sv:12:15
							localparam WORD_SIZE = _param_CC492_WORD_SIZE;
							// Trace: src/VX_cache_cluster.sv:13:15
							localparam CRSQ_SIZE = _param_CC492_CRSQ_SIZE;
							// Trace: src/VX_cache_cluster.sv:14:15
							localparam MSHR_SIZE = _param_CC492_MSHR_SIZE;
							// Trace: src/VX_cache_cluster.sv:15:15
							localparam MRSQ_SIZE = _param_CC492_MRSQ_SIZE;
							// Trace: src/VX_cache_cluster.sv:16:15
							localparam MREQ_SIZE = _param_CC492_MREQ_SIZE;
							// Trace: src/VX_cache_cluster.sv:17:15
							localparam WRITE_ENABLE = _param_CC492_WRITE_ENABLE;
							// Trace: src/VX_cache_cluster.sv:18:15
							localparam WRITEBACK = _param_CC492_WRITEBACK;
							// Trace: src/VX_cache_cluster.sv:19:15
							localparam DIRTY_BYTES = _param_CC492_DIRTY_BYTES;
							// Trace: src/VX_cache_cluster.sv:20:15
							localparam REPL_POLICY = _param_CC492_REPL_POLICY;
							// Trace: src/VX_cache_cluster.sv:21:15
							localparam VX_gpu_pkg_UUID_WIDTH = 1;
							localparam TAG_WIDTH = _param_CC492_TAG_WIDTH;
							// Trace: src/VX_cache_cluster.sv:22:15
							localparam NC_ENABLE = _param_CC492_NC_ENABLE;
							// Trace: src/VX_cache_cluster.sv:23:15
							localparam CORE_OUT_BUF = _param_CC492_CORE_OUT_BUF;
							// Trace: src/VX_cache_cluster.sv:24:15
							localparam MEM_OUT_BUF = _param_CC492_MEM_OUT_BUF;
							// Trace: src/VX_cache_cluster.sv:26:5
							wire clk;
							// Trace: src/VX_cache_cluster.sv:27:5
							wire reset;
							// Trace: src/VX_cache_cluster.sv:28:5
							localparam _mbase_core_bus_if = 0;
							// Trace: src/VX_cache_cluster.sv:29:5
							localparam _mbase_mem_bus_if = 0;
							// Trace: src/VX_cache_cluster.sv:31:5
							localparam NUM_CACHES = NUM_UNITS;
							// Trace: src/VX_cache_cluster.sv:32:5
							localparam PASSTHRU = 1'd0;
							// Trace: src/VX_cache_cluster.sv:33:5
							localparam ARB_TAG_WIDTH = 3;
							// Trace: src/VX_cache_cluster.sv:34:5
							localparam CACHE_MEM_TAG_WIDTH = 5;
							// Trace: src/VX_cache_cluster.sv:36:5
							localparam BYPASS_TAG_WIDTH = 5;
							// Trace: src/VX_cache_cluster.sv:38:5
							localparam NC_TAG_WIDTH = 6;
							// Trace: src/VX_cache_cluster.sv:39:5
							localparam MEM_TAG_WIDTH = (PASSTHRU ? BYPASS_TAG_WIDTH : (NC_ENABLE ? NC_TAG_WIDTH : CACHE_MEM_TAG_WIDTH));
							// Trace: src/VX_cache_cluster.sv:40:5
							// expanded interface instance: cache_mem_bus_if
							localparam _param_A4879_DATA_SIZE = LINE_SIZE;
							localparam _param_A4879_TAG_WIDTH = MEM_TAG_WIDTH;
							genvar _arr_A4879;
							for (_arr_A4879 = 0; _arr_A4879 <= 0; _arr_A4879 = _arr_A4879 + 1) begin : cache_mem_bus_if
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_A4879_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
								localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
								localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_A4879_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 26;
								// Trace: src/VX_mem_bus_if.sv:8:5
								localparam VX_gpu_pkg_UUID_WIDTH = 1;
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:12:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:20:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:24:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire [611:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire [517:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:30:5
								// Trace: src/VX_mem_bus_if.sv:38:5
							end
							// Trace: src/VX_cache_cluster.sv:44:5
							// expanded interface instance: arb_core_bus_if
							localparam _param_F9BC9_DATA_SIZE = WORD_SIZE;
							localparam _param_F9BC9_TAG_WIDTH = ARB_TAG_WIDTH;
							genvar _arr_F9BC9;
							for (_arr_F9BC9 = 0; _arr_F9BC9 <= 0; _arr_F9BC9 = _arr_F9BC9 + 1) begin : arb_core_bus_if
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_mem_bus_if.sv:2:15
								localparam DATA_SIZE = _param_F9BC9_DATA_SIZE;
								// Trace: src/VX_mem_bus_if.sv:3:15
								localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
								localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
								localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:4:15
								localparam TAG_WIDTH = _param_F9BC9_TAG_WIDTH;
								// Trace: src/VX_mem_bus_if.sv:5:15
								localparam MEM_ADDR_WIDTH = 32;
								// Trace: src/VX_mem_bus_if.sv:6:15
								localparam ADDR_WIDTH = 28;
								// Trace: src/VX_mem_bus_if.sv:8:5
								localparam VX_gpu_pkg_UUID_WIDTH = 1;
								// removed localparam type tag_t
								// Trace: src/VX_mem_bus_if.sv:12:5
								// removed localparam type req_data_t
								// Trace: src/VX_mem_bus_if.sv:20:5
								// removed localparam type rsp_data_t
								// Trace: src/VX_mem_bus_if.sv:24:5
								wire req_valid;
								// Trace: src/VX_mem_bus_if.sv:25:5
								wire [178:0] req_data;
								// Trace: src/VX_mem_bus_if.sv:26:5
								wire req_ready;
								// Trace: src/VX_mem_bus_if.sv:27:5
								wire rsp_valid;
								// Trace: src/VX_mem_bus_if.sv:28:5
								wire [130:0] rsp_data;
								// Trace: src/VX_mem_bus_if.sv:29:5
								wire rsp_ready;
								// Trace: src/VX_mem_bus_if.sv:30:5
								// Trace: src/VX_mem_bus_if.sv:38:5
							end
							// Trace: src/VX_cache_cluster.sv:48:5
							genvar _gv_i_191;
							for (_gv_i_191 = 0; _gv_i_191 < NUM_REQS; _gv_i_191 = _gv_i_191 + 1) begin : g_core_arb
								localparam i = _gv_i_191;
								// Trace: src/VX_cache_cluster.sv:49:9
								// expanded interface instance: core_bus_tmp_if
								localparam _param_A62F7_DATA_SIZE = WORD_SIZE;
								localparam _param_A62F7_TAG_WIDTH = TAG_WIDTH;
								genvar _arr_A62F7;
								for (_arr_A62F7 = 0; _arr_A62F7 <= 0; _arr_A62F7 = _arr_A62F7 + 1) begin : core_bus_tmp_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_A62F7_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_A62F7_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 28;
									// Trace: src/VX_mem_bus_if.sv:8:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:12:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:20:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:24:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire [178:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire [130:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:30:5
									// Trace: src/VX_mem_bus_if.sv:38:5
								end
								// Trace: src/VX_cache_cluster.sv:53:9
								// expanded interface instance: arb_core_bus_tmp_if
								localparam _param_E788B_DATA_SIZE = WORD_SIZE;
								localparam _param_E788B_TAG_WIDTH = ARB_TAG_WIDTH;
								genvar _arr_E788B;
								for (_arr_E788B = 0; _arr_E788B <= 0; _arr_E788B = _arr_E788B + 1) begin : arb_core_bus_tmp_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_E788B_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_E788B_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 28;
									// Trace: src/VX_mem_bus_if.sv:8:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:12:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:20:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:24:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire [178:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire [130:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:30:5
									// Trace: src/VX_mem_bus_if.sv:38:5
								end
								genvar _gv_j_19;
								for (_gv_j_19 = 0; _gv_j_19 < NUM_INPUTS; _gv_j_19 = _gv_j_19 + 1) begin : g_core_bus_tmp_if
									localparam j = _gv_j_19;
									// Trace: src/VX_cache_cluster.sv:58:5
									assign core_bus_tmp_if[j].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].req_valid;
									// Trace: src/VX_cache_cluster.sv:59:5
									assign core_bus_tmp_if[j].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].req_data;
									// Trace: src/VX_cache_cluster.sv:60:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].req_ready = core_bus_tmp_if[j].req_ready;
									// Trace: src/VX_cache_cluster.sv:61:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].rsp_valid = core_bus_tmp_if[j].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:62:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].rsp_data = core_bus_tmp_if[j].rsp_data;
									// Trace: src/VX_cache_cluster.sv:63:5
									assign core_bus_tmp_if[j].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((j * NUM_REQS) + i) + _mbase_core_bus_if].rsp_ready;
								end
								// Trace: src/VX_cache_cluster.sv:65:9
								// expanded module instance: core_arb
								localparam _bbase_856A9_bus_in_if = 0;
								localparam _bbase_856A9_bus_out_if = 0;
								localparam _param_856A9_NUM_INPUTS = NUM_INPUTS;
								localparam _param_856A9_NUM_OUTPUTS = NUM_CACHES;
								localparam _param_856A9_DATA_SIZE = WORD_SIZE;
								localparam _param_856A9_TAG_WIDTH = TAG_WIDTH;
								localparam _param_856A9_TAG_SEL_IDX = TAG_SEL_IDX;
								localparam _param_856A9_ARBITER = "R";
								localparam _param_856A9_REQ_OUT_BUF = 0;
								localparam _param_856A9_RSP_OUT_BUF = 0;
								if (1) begin : core_arb
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_arb.sv:2:15
									localparam NUM_INPUTS = _param_856A9_NUM_INPUTS;
									// Trace: src/VX_mem_arb.sv:3:15
									localparam NUM_OUTPUTS = _param_856A9_NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:4:15
									localparam DATA_SIZE = _param_856A9_DATA_SIZE;
									// Trace: src/VX_mem_arb.sv:5:15
									localparam TAG_WIDTH = _param_856A9_TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:6:15
									localparam TAG_SEL_IDX = _param_856A9_TAG_SEL_IDX;
									// Trace: src/VX_mem_arb.sv:7:15
									localparam REQ_OUT_BUF = _param_856A9_REQ_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:8:15
									localparam RSP_OUT_BUF = _param_856A9_RSP_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:9:15
									localparam ARBITER = _param_856A9_ARBITER;
									// Trace: src/VX_mem_arb.sv:10:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_arb.sv:11:15
									localparam ADDR_WIDTH = 28;
									// Trace: src/VX_mem_arb.sv:12:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_arb.sv:14:5
									wire clk;
									// Trace: src/VX_mem_arb.sv:15:5
									wire reset;
									// Trace: src/VX_mem_arb.sv:16:5
									localparam _mbase_bus_in_if = 0;
									// Trace: src/VX_mem_arb.sv:17:5
									localparam _mbase_bus_out_if = 0;
									// Trace: src/VX_mem_arb.sv:19:5
									localparam DATA_WIDTH = 128;
									// Trace: src/VX_mem_arb.sv:20:5
									localparam LOG_NUM_REQS = 0;
									// Trace: src/VX_mem_arb.sv:21:5
									localparam REQ_DATAW = 179;
									// Trace: src/VX_mem_arb.sv:22:5
									localparam RSP_DATAW = 131;
									// Trace: src/VX_mem_arb.sv:23:5
									localparam SEL_COUNT = NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:24:5
									wire [0:0] req_valid_in;
									// Trace: src/VX_mem_arb.sv:25:5
									wire [178:0] req_data_in;
									// Trace: src/VX_mem_arb.sv:26:5
									wire [0:0] req_ready_in;
									// Trace: src/VX_mem_arb.sv:27:5
									wire [0:0] req_valid_out;
									// Trace: src/VX_mem_arb.sv:28:5
									wire [178:0] req_data_out;
									// Trace: src/VX_mem_arb.sv:29:5
									wire [0:0] req_sel_out;
									// Trace: src/VX_mem_arb.sv:30:5
									wire [0:0] req_ready_out;
									// Trace: src/VX_mem_arb.sv:31:5
									genvar _gv_i_183;
									for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
										localparam i = _gv_i_183;
										// Trace: src/VX_mem_arb.sv:32:9
										assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].core_bus_tmp_if[i + _mbase_bus_in_if].req_valid;
										// Trace: src/VX_mem_arb.sv:33:9
										assign req_data_in[i * 179+:179] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].core_bus_tmp_if[i + _mbase_bus_in_if].req_data;
										// Trace: src/VX_mem_arb.sv:34:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].core_bus_tmp_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:36:5
									VX_stream_arb #(
										.NUM_INPUTS(NUM_INPUTS),
										.NUM_OUTPUTS(NUM_OUTPUTS),
										.DATAW(REQ_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(REQ_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(req_valid_in),
										.ready_in(req_ready_in),
										.data_in(req_data_in),
										.data_out(req_data_out),
										.sel_out(req_sel_out),
										.valid_out(req_valid_out),
										.ready_out(req_ready_out)
									);
									// Trace: src/VX_mem_arb.sv:53:5
									genvar _gv_i_184;
									for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
										localparam i = _gv_i_184;
										// Trace: src/VX_mem_arb.sv:54:9
										wire [2:0] req_tag_out;
										// Trace: src/VX_mem_arb.sv:55:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
										// Trace: src/VX_mem_arb.sv:56:9
										assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[178], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[177-:28], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[149-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[21-:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[5-:3], req_tag_out} = req_data_out[i * 179+:179];
										// Trace: src/VX_mem_arb.sv:64:9
										assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
										if (1) begin : g_req_tag_out
											// Trace: src/VX_mem_arb.sv:76:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].req_data[2-:3] = req_tag_out;
										end
									end
									// Trace: src/VX_mem_arb.sv:79:5
									wire [0:0] rsp_valid_out;
									// Trace: src/VX_mem_arb.sv:80:5
									wire [130:0] rsp_data_out;
									// Trace: src/VX_mem_arb.sv:81:5
									wire [0:0] rsp_ready_out;
									// Trace: src/VX_mem_arb.sv:82:5
									wire [0:0] rsp_valid_in;
									// Trace: src/VX_mem_arb.sv:83:5
									wire [130:0] rsp_data_in;
									// Trace: src/VX_mem_arb.sv:84:5
									wire [0:0] rsp_ready_in;
									// Trace: src/VX_mem_arb.sv:85:5
									if (1) begin : g_rsp_arb
										genvar _gv_i_186;
										for (_gv_i_186 = 0; _gv_i_186 < NUM_OUTPUTS; _gv_i_186 = _gv_i_186 + 1) begin : g_rsp_data_in
											localparam i = _gv_i_186;
											// Trace: src/VX_mem_arb.sv:120:13
											assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
											// Trace: src/VX_mem_arb.sv:121:13
											assign rsp_data_in[i * 131+:131] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
											// Trace: src/VX_mem_arb.sv:122:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].arb_core_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
										end
										// Trace: src/VX_mem_arb.sv:124:9
										VX_stream_arb #(
											.NUM_INPUTS(NUM_OUTPUTS),
											.NUM_OUTPUTS(NUM_INPUTS),
											.DATAW(RSP_DATAW),
											.ARBITER(ARBITER),
											.OUT_BUF(RSP_OUT_BUF)
										) req_arb(
											.clk(clk),
											.reset(reset),
											.valid_in(rsp_valid_in),
											.ready_in(rsp_ready_in),
											.data_in(rsp_data_in),
											.data_out(rsp_data_out),
											.valid_out(rsp_valid_out),
											.ready_out(rsp_ready_out),
											.sel_out()
										);
									end
									// Trace: src/VX_mem_arb.sv:142:5
									genvar _gv_i_187;
									for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
										localparam i = _gv_i_187;
										// Trace: src/VX_mem_arb.sv:143:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].core_bus_tmp_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
										// Trace: src/VX_mem_arb.sv:144:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].core_bus_tmp_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 131+:131];
										// Trace: src/VX_mem_arb.sv:145:9
										assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_core_arb[_gv_i_191].core_bus_tmp_if[i + _mbase_bus_in_if].rsp_ready;
									end
								end
								assign core_arb.clk = clk;
								assign core_arb.reset = reset;
								genvar _gv_k_1;
								for (_gv_k_1 = 0; _gv_k_1 < NUM_CACHES; _gv_k_1 = _gv_k_1 + 1) begin : g_arb_core_bus_if
									localparam k = _gv_k_1;
									// Trace: src/VX_cache_cluster.sv:81:5
									assign arb_core_bus_if[(k * NUM_REQS) + i].req_valid = arb_core_bus_tmp_if[k].req_valid;
									// Trace: src/VX_cache_cluster.sv:82:5
									assign arb_core_bus_if[(k * NUM_REQS) + i].req_data = arb_core_bus_tmp_if[k].req_data;
									// Trace: src/VX_cache_cluster.sv:83:5
									assign arb_core_bus_tmp_if[k].req_ready = arb_core_bus_if[(k * NUM_REQS) + i].req_ready;
									// Trace: src/VX_cache_cluster.sv:84:5
									assign arb_core_bus_tmp_if[k].rsp_valid = arb_core_bus_if[(k * NUM_REQS) + i].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:85:5
									assign arb_core_bus_tmp_if[k].rsp_data = arb_core_bus_if[(k * NUM_REQS) + i].rsp_data;
									// Trace: src/VX_cache_cluster.sv:86:5
									assign arb_core_bus_if[(k * NUM_REQS) + i].rsp_ready = arb_core_bus_tmp_if[k].rsp_ready;
								end
							end
							// Trace: src/VX_cache_cluster.sv:89:6
							genvar _gv_i_192;
							for (_gv_i_192 = 0; _gv_i_192 < NUM_CACHES; _gv_i_192 = _gv_i_192 + 1) begin : g_cache_wrap
								localparam i = _gv_i_192;
								// Trace: src/VX_cache_cluster.sv:90:9
								// expanded module instance: cache_wrap
								localparam _bbase_665FE_core_bus_if = i * NUM_REQS;
								localparam _bbase_665FE_mem_bus_if = i * MEM_PORTS;
								localparam _param_665FE_INSTANCE_ID = "";
								localparam _param_665FE_CACHE_SIZE = CACHE_SIZE;
								localparam _param_665FE_LINE_SIZE = LINE_SIZE;
								localparam _param_665FE_NUM_BANKS = NUM_BANKS;
								localparam _param_665FE_NUM_WAYS = NUM_WAYS;
								localparam _param_665FE_WORD_SIZE = WORD_SIZE;
								localparam _param_665FE_NUM_REQS = NUM_REQS;
								localparam _param_665FE_MEM_PORTS = MEM_PORTS;
								localparam _param_665FE_WRITE_ENABLE = WRITE_ENABLE;
								localparam _param_665FE_WRITEBACK = WRITEBACK;
								localparam _param_665FE_DIRTY_BYTES = DIRTY_BYTES;
								localparam _param_665FE_REPL_POLICY = REPL_POLICY;
								localparam _param_665FE_CRSQ_SIZE = CRSQ_SIZE;
								localparam _param_665FE_MSHR_SIZE = MSHR_SIZE;
								localparam _param_665FE_MRSQ_SIZE = MRSQ_SIZE;
								localparam _param_665FE_MREQ_SIZE = MREQ_SIZE;
								localparam _param_665FE_TAG_WIDTH = ARB_TAG_WIDTH;
								localparam _param_665FE_TAG_SEL_IDX = TAG_SEL_IDX;
								localparam _param_665FE_CORE_OUT_BUF = CORE_OUT_BUF;
								localparam _param_665FE_MEM_OUT_BUF = MEM_OUT_BUF;
								localparam _param_665FE_NC_ENABLE = NC_ENABLE;
								localparam _param_665FE_PASSTHRU = PASSTHRU;
								if (1) begin : cache_wrap
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_cache_wrap.sv:2:15
									localparam INSTANCE_ID = _param_665FE_INSTANCE_ID;
									// Trace: src/VX_cache_wrap.sv:3:15
									localparam TAG_SEL_IDX = _param_665FE_TAG_SEL_IDX;
									// Trace: src/VX_cache_wrap.sv:4:15
									localparam NUM_REQS = _param_665FE_NUM_REQS;
									// Trace: src/VX_cache_wrap.sv:5:15
									localparam MEM_PORTS = _param_665FE_MEM_PORTS;
									// Trace: src/VX_cache_wrap.sv:6:15
									localparam CACHE_SIZE = _param_665FE_CACHE_SIZE;
									// Trace: src/VX_cache_wrap.sv:7:15
									localparam LINE_SIZE = _param_665FE_LINE_SIZE;
									// Trace: src/VX_cache_wrap.sv:8:15
									localparam NUM_BANKS = _param_665FE_NUM_BANKS;
									// Trace: src/VX_cache_wrap.sv:9:15
									localparam NUM_WAYS = _param_665FE_NUM_WAYS;
									// Trace: src/VX_cache_wrap.sv:10:15
									localparam WORD_SIZE = _param_665FE_WORD_SIZE;
									// Trace: src/VX_cache_wrap.sv:11:15
									localparam CRSQ_SIZE = _param_665FE_CRSQ_SIZE;
									// Trace: src/VX_cache_wrap.sv:12:15
									localparam MSHR_SIZE = _param_665FE_MSHR_SIZE;
									// Trace: src/VX_cache_wrap.sv:13:15
									localparam MRSQ_SIZE = _param_665FE_MRSQ_SIZE;
									// Trace: src/VX_cache_wrap.sv:14:15
									localparam MREQ_SIZE = _param_665FE_MREQ_SIZE;
									// Trace: src/VX_cache_wrap.sv:15:15
									localparam WRITE_ENABLE = _param_665FE_WRITE_ENABLE;
									// Trace: src/VX_cache_wrap.sv:16:15
									localparam WRITEBACK = _param_665FE_WRITEBACK;
									// Trace: src/VX_cache_wrap.sv:17:15
									localparam DIRTY_BYTES = _param_665FE_DIRTY_BYTES;
									// Trace: src/VX_cache_wrap.sv:18:15
									localparam REPL_POLICY = _param_665FE_REPL_POLICY;
									// Trace: src/VX_cache_wrap.sv:19:15
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									localparam TAG_WIDTH = _param_665FE_TAG_WIDTH;
									// Trace: src/VX_cache_wrap.sv:20:15
									localparam NC_ENABLE = _param_665FE_NC_ENABLE;
									// Trace: src/VX_cache_wrap.sv:21:15
									localparam PASSTHRU = _param_665FE_PASSTHRU;
									// Trace: src/VX_cache_wrap.sv:22:15
									localparam CORE_OUT_BUF = _param_665FE_CORE_OUT_BUF;
									// Trace: src/VX_cache_wrap.sv:23:15
									localparam MEM_OUT_BUF = _param_665FE_MEM_OUT_BUF;
									// Trace: src/VX_cache_wrap.sv:25:5
									wire clk;
									// Trace: src/VX_cache_wrap.sv:26:5
									wire reset;
									// Trace: src/VX_cache_wrap.sv:27:5
									localparam _mbase_core_bus_if = _bbase_665FE_core_bus_if;
									// Trace: src/VX_cache_wrap.sv:28:5
									localparam _mbase_mem_bus_if = _bbase_665FE_mem_bus_if;
									// Trace: src/VX_cache_wrap.sv:30:5
									localparam CACHE_MEM_TAG_WIDTH = 5;
									// Trace: src/VX_cache_wrap.sv:32:5
									localparam BYPASS_TAG_WIDTH = 5;
									// Trace: src/VX_cache_wrap.sv:34:5
									localparam NC_TAG_WIDTH = 6;
									// Trace: src/VX_cache_wrap.sv:35:5
									localparam MEM_TAG_WIDTH = (PASSTHRU ? BYPASS_TAG_WIDTH : (NC_ENABLE ? NC_TAG_WIDTH : CACHE_MEM_TAG_WIDTH));
									// Trace: src/VX_cache_wrap.sv:36:5
									localparam BYPASS_ENABLE = 1'd1;
									// Trace: src/VX_cache_wrap.sv:37:5
									// expanded interface instance: core_bus_cache_if
									localparam _param_24C1C_DATA_SIZE = WORD_SIZE;
									localparam _param_24C1C_TAG_WIDTH = TAG_WIDTH;
									genvar _arr_24C1C;
									for (_arr_24C1C = 0; _arr_24C1C <= 0; _arr_24C1C = _arr_24C1C + 1) begin : core_bus_cache_if
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_24C1C_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_24C1C_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 28;
										// Trace: src/VX_mem_bus_if.sv:8:5
										localparam VX_gpu_pkg_UUID_WIDTH = 1;
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:12:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:20:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:24:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire [178:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire [130:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:30:5
										// Trace: src/VX_mem_bus_if.sv:38:5
									end
									// Trace: src/VX_cache_wrap.sv:41:5
									// expanded interface instance: mem_bus_cache_if
									localparam _param_D895D_DATA_SIZE = LINE_SIZE;
									localparam _param_D895D_TAG_WIDTH = CACHE_MEM_TAG_WIDTH;
									genvar _arr_D895D;
									for (_arr_D895D = 0; _arr_D895D <= 0; _arr_D895D = _arr_D895D + 1) begin : mem_bus_cache_if
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_D895D_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_D895D_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 26;
										// Trace: src/VX_mem_bus_if.sv:8:5
										localparam VX_gpu_pkg_UUID_WIDTH = 1;
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:12:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:20:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:24:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire [610:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire [516:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:30:5
										// Trace: src/VX_mem_bus_if.sv:38:5
									end
									// Trace: src/VX_cache_wrap.sv:45:5
									// expanded interface instance: mem_bus_tmp_if
									localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
									localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH;
									genvar _arr_4FE36;
									for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 26;
										// Trace: src/VX_mem_bus_if.sv:8:5
										localparam VX_gpu_pkg_UUID_WIDTH = 1;
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:12:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:20:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:24:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire [611:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire [517:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:30:5
										// Trace: src/VX_mem_bus_if.sv:38:5
									end
									// Trace: src/VX_cache_wrap.sv:49:5
									if (BYPASS_ENABLE) begin : g_bypass
										// Trace: src/VX_cache_wrap.sv:50:9
										// expanded module instance: cache_bypass
										localparam _bbase_714AA_core_bus_in_if = i * NUM_REQS;
										localparam _bbase_714AA_core_bus_out_if = 0;
										localparam _bbase_714AA_mem_bus_in_if = 0;
										localparam _bbase_714AA_mem_bus_out_if = 0;
										localparam _param_714AA_NUM_REQS = NUM_REQS;
										localparam _param_714AA_MEM_PORTS = MEM_PORTS;
										localparam _param_714AA_TAG_SEL_IDX = TAG_SEL_IDX;
										localparam _param_714AA_CACHE_ENABLE = !PASSTHRU;
										localparam _param_714AA_WORD_SIZE = WORD_SIZE;
										localparam _param_714AA_LINE_SIZE = LINE_SIZE;
										localparam _param_714AA_CORE_ADDR_WIDTH = 28;
										localparam _param_714AA_CORE_TAG_WIDTH = TAG_WIDTH;
										localparam _param_714AA_MEM_ADDR_WIDTH = 26;
										localparam _param_714AA_MEM_TAG_IN_WIDTH = CACHE_MEM_TAG_WIDTH;
										localparam _param_714AA_CORE_OUT_BUF = CORE_OUT_BUF;
										localparam _param_714AA_MEM_OUT_BUF = MEM_OUT_BUF;
										if (1) begin : cache_bypass
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_cache_bypass.sv:2:15
											localparam NUM_REQS = _param_714AA_NUM_REQS;
											// Trace: src/VX_cache_bypass.sv:3:15
											localparam MEM_PORTS = _param_714AA_MEM_PORTS;
											// Trace: src/VX_cache_bypass.sv:4:15
											localparam TAG_SEL_IDX = _param_714AA_TAG_SEL_IDX;
											// Trace: src/VX_cache_bypass.sv:5:15
											localparam CACHE_ENABLE = _param_714AA_CACHE_ENABLE;
											// Trace: src/VX_cache_bypass.sv:6:15
											localparam WORD_SIZE = _param_714AA_WORD_SIZE;
											// Trace: src/VX_cache_bypass.sv:7:15
											localparam LINE_SIZE = _param_714AA_LINE_SIZE;
											// Trace: src/VX_cache_bypass.sv:8:15
											localparam CORE_ADDR_WIDTH = _param_714AA_CORE_ADDR_WIDTH;
											// Trace: src/VX_cache_bypass.sv:9:15
											localparam CORE_TAG_WIDTH = _param_714AA_CORE_TAG_WIDTH;
											// Trace: src/VX_cache_bypass.sv:10:15
											localparam MEM_ADDR_WIDTH = _param_714AA_MEM_ADDR_WIDTH;
											// Trace: src/VX_cache_bypass.sv:11:15
											localparam MEM_TAG_IN_WIDTH = _param_714AA_MEM_TAG_IN_WIDTH;
											// Trace: src/VX_cache_bypass.sv:12:15
											localparam CORE_OUT_BUF = _param_714AA_CORE_OUT_BUF;
											// Trace: src/VX_cache_bypass.sv:13:15
											localparam MEM_OUT_BUF = _param_714AA_MEM_OUT_BUF;
											// Trace: src/VX_cache_bypass.sv:15:5
											wire clk;
											// Trace: src/VX_cache_bypass.sv:16:5
											wire reset;
											// Trace: src/VX_cache_bypass.sv:17:5
											localparam _mbase_core_bus_in_if = _bbase_714AA_core_bus_in_if;
											// Trace: src/VX_cache_bypass.sv:18:5
											localparam _mbase_core_bus_out_if = 0;
											// Trace: src/VX_cache_bypass.sv:19:5
											localparam _mbase_mem_bus_in_if = 0;
											// Trace: src/VX_cache_bypass.sv:20:5
											localparam _mbase_mem_bus_out_if = 0;
											// Trace: src/VX_cache_bypass.sv:22:5
											localparam DIRECT_PASSTHRU = (!CACHE_ENABLE && 1'd0) && 1'd1;
											// Trace: src/VX_cache_bypass.sv:23:5
											localparam CORE_DATA_WIDTH = 128;
											// Trace: src/VX_cache_bypass.sv:24:5
											localparam WORDS_PER_LINE = 4;
											// Trace: src/VX_cache_bypass.sv:25:5
											localparam WSEL_BITS = 2;
											// Trace: src/VX_cache_bypass.sv:26:5
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam CORE_TAG_ID_WIDTH = 2;
											// Trace: src/VX_cache_bypass.sv:27:5
											localparam MEM_TAG_ID_WIDTH = 2;
											// Trace: src/VX_cache_bypass.sv:28:5
											localparam MEM_TAG_NC1_WIDTH = 3;
											// Trace: src/VX_cache_bypass.sv:29:5
											localparam MEM_TAG_NC2_WIDTH = 5;
											// Trace: src/VX_cache_bypass.sv:30:5
											localparam MEM_TAG_OUT_WIDTH = (CACHE_ENABLE ? MEM_TAG_NC2_WIDTH : MEM_TAG_NC2_WIDTH);
											// Trace: src/VX_cache_bypass.sv:31:5
											// expanded interface instance: core_bus_nc_switch_if
											localparam _param_95306_DATA_SIZE = WORD_SIZE;
											localparam _param_95306_TAG_WIDTH = CORE_TAG_WIDTH;
											genvar _arr_95306;
											for (_arr_95306 = 0; _arr_95306 <= (((CACHE_ENABLE ? 2 : 1) * NUM_REQS) - 1); _arr_95306 = _arr_95306 + 1) begin : core_bus_nc_switch_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_95306_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_95306_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 28;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [178:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [130:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache_bypass.sv:35:5
											wire [0:0] core_req_nc_sel;
											// Trace: src/VX_cache_bypass.sv:36:5
											genvar _gv_i_56;
											localparam VX_gpu_pkg_MEM_REQ_FLAG_IO = 1;
											for (_gv_i_56 = 0; _gv_i_56 < NUM_REQS; _gv_i_56 = _gv_i_56 + 1) begin : g_core_req_is_nc
												localparam i = _gv_i_56;
												if (CACHE_ENABLE) begin : g_cache
													// Trace: src/VX_cache_bypass.sv:38:13
													assign core_req_nc_sel[i] = ~Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_in_if].req_data[4];
												end
												else begin : g_no_cache
													// Trace: src/VX_cache_bypass.sv:40:13
													assign core_req_nc_sel[i] = 1'b0;
												end
											end
											// Trace: src/VX_cache_bypass.sv:43:5
											// expanded module instance: core_bus_nc_switch
											localparam _bbase_69FDB_bus_in_if = i * NUM_REQS;
											localparam _bbase_69FDB_bus_out_if = 0;
											localparam _param_69FDB_NUM_INPUTS = NUM_REQS;
											localparam _param_69FDB_NUM_OUTPUTS = (CACHE_ENABLE ? 2 : 1) * NUM_REQS;
											localparam _param_69FDB_DATA_SIZE = WORD_SIZE;
											localparam _param_69FDB_TAG_WIDTH = CORE_TAG_WIDTH;
											localparam _param_69FDB_ARBITER = "R";
											localparam _param_69FDB_REQ_OUT_BUF = 0;
											localparam _param_69FDB_RSP_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
											if (1) begin : core_bus_nc_switch
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_switch.sv:2:15
												localparam NUM_INPUTS = _param_69FDB_NUM_INPUTS;
												// Trace: src/VX_mem_switch.sv:3:15
												localparam NUM_OUTPUTS = _param_69FDB_NUM_OUTPUTS;
												// Trace: src/VX_mem_switch.sv:4:15
												localparam DATA_SIZE = _param_69FDB_DATA_SIZE;
												// Trace: src/VX_mem_switch.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_switch.sv:6:15
												localparam ADDR_WIDTH = 28;
												// Trace: src/VX_mem_switch.sv:7:15
												localparam TAG_WIDTH = _param_69FDB_TAG_WIDTH;
												// Trace: src/VX_mem_switch.sv:8:15
												localparam REQ_OUT_BUF = _param_69FDB_REQ_OUT_BUF;
												// Trace: src/VX_mem_switch.sv:9:15
												localparam RSP_OUT_BUF = _param_69FDB_RSP_OUT_BUF;
												// Trace: src/VX_mem_switch.sv:10:15
												localparam ARBITER = _param_69FDB_ARBITER;
												// Trace: src/VX_mem_switch.sv:11:15
												localparam NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? ((NUM_INPUTS + NUM_OUTPUTS) - 1) / NUM_OUTPUTS : ((NUM_OUTPUTS + NUM_INPUTS) - 1) / NUM_INPUTS);
												// Trace: src/VX_mem_switch.sv:12:15
												localparam SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
												// Trace: src/VX_mem_switch.sv:13:15
												localparam LOG_NUM_REQS = $clog2(NUM_REQS);
												// Trace: src/VX_mem_switch.sv:15:5
												wire clk;
												// Trace: src/VX_mem_switch.sv:16:5
												wire reset;
												// Trace: src/VX_mem_switch.sv:17:5
												wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] bus_sel;
												// Trace: src/VX_mem_switch.sv:18:5
												localparam _mbase_bus_in_if = _bbase_69FDB_bus_in_if;
												// Trace: src/VX_mem_switch.sv:19:5
												localparam _mbase_bus_out_if = 0;
												// Trace: src/VX_mem_switch.sv:21:5
												localparam DATA_WIDTH = 128;
												// Trace: src/VX_mem_switch.sv:22:5
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam REQ_DATAW = 179;
												// Trace: src/VX_mem_switch.sv:23:5
												localparam RSP_DATAW = 131;
												// Trace: src/VX_mem_switch.sv:24:5
												wire [0:0] req_valid_in;
												// Trace: src/VX_mem_switch.sv:25:5
												wire [178:0] req_data_in;
												// Trace: src/VX_mem_switch.sv:26:5
												wire [0:0] req_ready_in;
												// Trace: src/VX_mem_switch.sv:27:5
												wire [NUM_OUTPUTS - 1:0] req_valid_out;
												// Trace: src/VX_mem_switch.sv:28:5
												wire [(NUM_OUTPUTS * 179) - 1:0] req_data_out;
												// Trace: src/VX_mem_switch.sv:29:5
												wire [NUM_OUTPUTS - 1:0] req_ready_out;
												// Trace: src/VX_mem_switch.sv:30:5
												genvar _gv_i_109;
												for (_gv_i_109 = 0; _gv_i_109 < NUM_INPUTS; _gv_i_109 = _gv_i_109 + 1) begin : g_req_data_in
													localparam i = _gv_i_109;
													// Trace: src/VX_mem_switch.sv:31:9
													assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_bus_in_if].req_valid;
													// Trace: src/VX_mem_switch.sv:32:9
													assign req_data_in[i * 179+:179] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_bus_in_if].req_data;
													// Trace: src/VX_mem_switch.sv:33:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
												end
												// Trace: src/VX_mem_switch.sv:35:5
												VX_stream_switch #(
													.NUM_INPUTS(NUM_INPUTS),
													.NUM_OUTPUTS(NUM_OUTPUTS),
													.DATAW(REQ_DATAW),
													.OUT_BUF(REQ_OUT_BUF)
												) req_switch(
													.clk(clk),
													.reset(reset),
													.sel_in(bus_sel),
													.valid_in(req_valid_in),
													.data_in(req_data_in),
													.ready_in(req_ready_in),
													.valid_out(req_valid_out),
													.data_out(req_data_out),
													.ready_out(req_ready_out)
												);
												// Trace: src/VX_mem_switch.sv:51:5
												genvar _gv_i_110;
												for (_gv_i_110 = 0; _gv_i_110 < NUM_OUTPUTS; _gv_i_110 = _gv_i_110 + 1) begin : g_req_data_out
													localparam i = _gv_i_110;
													// Trace: src/VX_mem_switch.sv:52:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
													// Trace: src/VX_mem_switch.sv:53:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_data = req_data_out[i * 179+:179];
													// Trace: src/VX_mem_switch.sv:54:9
													assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].req_ready;
												end
												// Trace: src/VX_mem_switch.sv:56:5
												wire [NUM_OUTPUTS - 1:0] rsp_valid_in;
												// Trace: src/VX_mem_switch.sv:57:5
												wire [(NUM_OUTPUTS * 131) - 1:0] rsp_data_in;
												// Trace: src/VX_mem_switch.sv:58:5
												wire [NUM_OUTPUTS - 1:0] rsp_ready_in;
												// Trace: src/VX_mem_switch.sv:59:5
												wire [0:0] rsp_valid_out;
												// Trace: src/VX_mem_switch.sv:60:5
												wire [130:0] rsp_data_out;
												// Trace: src/VX_mem_switch.sv:61:5
												wire [0:0] rsp_ready_out;
												// Trace: src/VX_mem_switch.sv:62:5
												genvar _gv_i_111;
												for (_gv_i_111 = 0; _gv_i_111 < NUM_OUTPUTS; _gv_i_111 = _gv_i_111 + 1) begin : g_rsp_data_in
													localparam i = _gv_i_111;
													// Trace: src/VX_mem_switch.sv:63:9
													assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_valid;
													// Trace: src/VX_mem_switch.sv:64:9
													assign rsp_data_in[i * 131+:131] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_data;
													// Trace: src/VX_mem_switch.sv:65:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_switch_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
												end
												// Trace: src/VX_mem_switch.sv:67:5
												VX_stream_arb #(
													.NUM_INPUTS(NUM_OUTPUTS),
													.NUM_OUTPUTS(NUM_INPUTS),
													.DATAW(RSP_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(RSP_OUT_BUF)
												) rsp_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(rsp_valid_in),
													.data_in(rsp_data_in),
													.ready_in(rsp_ready_in),
													.valid_out(rsp_valid_out),
													.data_out(rsp_data_out),
													.ready_out(rsp_ready_out),
													.sel_out()
												);
												// Trace: src/VX_mem_switch.sv:84:5
												genvar _gv_i_112;
												for (_gv_i_112 = 0; _gv_i_112 < NUM_INPUTS; _gv_i_112 = _gv_i_112 + 1) begin : g_rsp_data_out
													localparam i = _gv_i_112;
													// Trace: src/VX_mem_switch.sv:85:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
													// Trace: src/VX_mem_switch.sv:86:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 131+:131];
													// Trace: src/VX_mem_switch.sv:87:9
													assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_bus_in_if].rsp_ready;
												end
											end
											assign core_bus_nc_switch.clk = clk;
											assign core_bus_nc_switch.reset = reset;
											assign core_bus_nc_switch.bus_sel = core_req_nc_sel;
											// Trace: src/VX_cache_bypass.sv:58:5
											// expanded interface instance: core_bus_in_nc_if
											localparam _param_C0263_DATA_SIZE = WORD_SIZE;
											localparam _param_C0263_TAG_WIDTH = CORE_TAG_WIDTH;
											genvar _arr_C0263;
											for (_arr_C0263 = 0; _arr_C0263 <= 0; _arr_C0263 = _arr_C0263 + 1) begin : core_bus_in_nc_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_C0263_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_C0263_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 28;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [178:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [130:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache_bypass.sv:62:5
											genvar _gv_i_57;
											for (_gv_i_57 = 0; _gv_i_57 < NUM_REQS; _gv_i_57 = _gv_i_57 + 1) begin : g_core_bus_nc_switch_if
												localparam i = _gv_i_57;
												// Trace: src/VX_cache_bypass.sv:63:9
												assign core_bus_in_nc_if[i].req_valid = core_bus_nc_switch_if[0 + i].req_valid;
												// Trace: src/VX_cache_bypass.sv:64:9
												assign core_bus_in_nc_if[i].req_data = core_bus_nc_switch_if[0 + i].req_data;
												// Trace: src/VX_cache_bypass.sv:65:9
												assign core_bus_nc_switch_if[0 + i].req_ready = core_bus_in_nc_if[i].req_ready;
												// Trace: src/VX_cache_bypass.sv:66:9
												assign core_bus_nc_switch_if[0 + i].rsp_valid = core_bus_in_nc_if[i].rsp_valid;
												// Trace: src/VX_cache_bypass.sv:67:9
												assign core_bus_nc_switch_if[0 + i].rsp_data = core_bus_in_nc_if[i].rsp_data;
												// Trace: src/VX_cache_bypass.sv:68:9
												assign core_bus_in_nc_if[i].rsp_ready = core_bus_nc_switch_if[0 + i].rsp_ready;
												if (CACHE_ENABLE) begin : g_cache
													// Trace: src/VX_cache_bypass.sv:70:13
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = core_bus_nc_switch_if[1 + i].req_valid;
													// Trace: src/VX_cache_bypass.sv:71:13
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = core_bus_nc_switch_if[1 + i].req_data;
													// Trace: src/VX_cache_bypass.sv:72:13
													assign core_bus_nc_switch_if[1 + i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_ready;
													// Trace: src/VX_cache_bypass.sv:73:13
													assign core_bus_nc_switch_if[1 + i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_valid;
													// Trace: src/VX_cache_bypass.sv:74:13
													assign core_bus_nc_switch_if[1 + i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_data;
													// Trace: src/VX_cache_bypass.sv:75:13
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = core_bus_nc_switch_if[1 + i].rsp_ready;
												end
												else begin : g_no_cache
													// Trace: src/VX_cache_bypass.sv:77:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_valid = 0;
													// Trace: src/VX_cache_bypass.sv:78:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].req_data = 1'sb0;
													// Trace: src/VX_cache_bypass.sv:79:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_out_if].rsp_ready = 0;
												end
											end
											// Trace: src/VX_cache_bypass.sv:82:5
											// expanded interface instance: core_bus_nc_arb_if
											localparam _param_D50AC_DATA_SIZE = WORD_SIZE;
											localparam _param_D50AC_TAG_WIDTH = MEM_TAG_NC1_WIDTH;
											genvar _arr_D50AC;
											for (_arr_D50AC = 0; _arr_D50AC <= 0; _arr_D50AC = _arr_D50AC + 1) begin : core_bus_nc_arb_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_D50AC_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_D50AC_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 28;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [178:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [130:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache_bypass.sv:86:5
											// expanded module instance: core_bus_nc_arb
											localparam _bbase_1376F_bus_in_if = 0;
											localparam _bbase_1376F_bus_out_if = 0;
											localparam _param_1376F_NUM_INPUTS = NUM_REQS;
											localparam _param_1376F_NUM_OUTPUTS = MEM_PORTS;
											localparam _param_1376F_DATA_SIZE = WORD_SIZE;
											localparam _param_1376F_TAG_WIDTH = CORE_TAG_WIDTH;
											localparam _param_1376F_TAG_SEL_IDX = TAG_SEL_IDX;
											localparam _param_1376F_ARBITER = (CACHE_ENABLE ? "P" : "R");
											localparam _param_1376F_REQ_OUT_BUF = 0;
											localparam _param_1376F_RSP_OUT_BUF = 0;
											if (1) begin : core_bus_nc_arb
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_arb.sv:2:15
												localparam NUM_INPUTS = _param_1376F_NUM_INPUTS;
												// Trace: src/VX_mem_arb.sv:3:15
												localparam NUM_OUTPUTS = _param_1376F_NUM_OUTPUTS;
												// Trace: src/VX_mem_arb.sv:4:15
												localparam DATA_SIZE = _param_1376F_DATA_SIZE;
												// Trace: src/VX_mem_arb.sv:5:15
												localparam TAG_WIDTH = _param_1376F_TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:6:15
												localparam TAG_SEL_IDX = _param_1376F_TAG_SEL_IDX;
												// Trace: src/VX_mem_arb.sv:7:15
												localparam REQ_OUT_BUF = _param_1376F_REQ_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:8:15
												localparam RSP_OUT_BUF = _param_1376F_RSP_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:9:15
												localparam ARBITER = _param_1376F_ARBITER;
												// Trace: src/VX_mem_arb.sv:10:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_arb.sv:11:15
												localparam ADDR_WIDTH = 28;
												// Trace: src/VX_mem_arb.sv:12:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_arb.sv:14:5
												wire clk;
												// Trace: src/VX_mem_arb.sv:15:5
												wire reset;
												// Trace: src/VX_mem_arb.sv:16:5
												localparam _mbase_bus_in_if = 0;
												// Trace: src/VX_mem_arb.sv:17:5
												localparam _mbase_bus_out_if = 0;
												// Trace: src/VX_mem_arb.sv:19:5
												localparam DATA_WIDTH = 128;
												// Trace: src/VX_mem_arb.sv:20:5
												localparam LOG_NUM_REQS = 0;
												// Trace: src/VX_mem_arb.sv:21:5
												localparam REQ_DATAW = 179;
												// Trace: src/VX_mem_arb.sv:22:5
												localparam RSP_DATAW = 131;
												// Trace: src/VX_mem_arb.sv:23:5
												localparam SEL_COUNT = NUM_OUTPUTS;
												// Trace: src/VX_mem_arb.sv:24:5
												wire [0:0] req_valid_in;
												// Trace: src/VX_mem_arb.sv:25:5
												wire [178:0] req_data_in;
												// Trace: src/VX_mem_arb.sv:26:5
												wire [0:0] req_ready_in;
												// Trace: src/VX_mem_arb.sv:27:5
												wire [0:0] req_valid_out;
												// Trace: src/VX_mem_arb.sv:28:5
												wire [178:0] req_data_out;
												// Trace: src/VX_mem_arb.sv:29:5
												wire [0:0] req_sel_out;
												// Trace: src/VX_mem_arb.sv:30:5
												wire [0:0] req_ready_out;
												// Trace: src/VX_mem_arb.sv:31:5
												genvar _gv_i_183;
												for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
													localparam i = _gv_i_183;
													// Trace: src/VX_mem_arb.sv:32:9
													assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_valid;
													// Trace: src/VX_mem_arb.sv:33:9
													assign req_data_in[i * 179+:179] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_data;
													// Trace: src/VX_mem_arb.sv:34:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
												end
												// Trace: src/VX_mem_arb.sv:36:5
												VX_stream_arb #(
													.NUM_INPUTS(NUM_INPUTS),
													.NUM_OUTPUTS(NUM_OUTPUTS),
													.DATAW(REQ_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(REQ_OUT_BUF)
												) req_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(req_valid_in),
													.ready_in(req_ready_in),
													.data_in(req_data_in),
													.data_out(req_data_out),
													.sel_out(req_sel_out),
													.valid_out(req_valid_out),
													.ready_out(req_ready_out)
												);
												// Trace: src/VX_mem_arb.sv:53:5
												genvar _gv_i_184;
												for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
													localparam i = _gv_i_184;
													// Trace: src/VX_mem_arb.sv:54:9
													wire [2:0] req_tag_out;
													// Trace: src/VX_mem_arb.sv:55:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
													// Trace: src/VX_mem_arb.sv:56:9
													assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[178], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[177-:28], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[149-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[21-:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[5-:3], req_tag_out} = req_data_out[i * 179+:179];
													// Trace: src/VX_mem_arb.sv:64:9
													assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_ready;
													if (1) begin : g_req_tag_out
														// Trace: src/VX_mem_arb.sv:76:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].req_data[2-:3] = req_tag_out;
													end
												end
												// Trace: src/VX_mem_arb.sv:79:5
												wire [0:0] rsp_valid_out;
												// Trace: src/VX_mem_arb.sv:80:5
												wire [130:0] rsp_data_out;
												// Trace: src/VX_mem_arb.sv:81:5
												wire [0:0] rsp_ready_out;
												// Trace: src/VX_mem_arb.sv:82:5
												wire [0:0] rsp_valid_in;
												// Trace: src/VX_mem_arb.sv:83:5
												wire [130:0] rsp_data_in;
												// Trace: src/VX_mem_arb.sv:84:5
												wire [0:0] rsp_ready_in;
												// Trace: src/VX_mem_arb.sv:85:5
												if (1) begin : g_rsp_arb
													genvar _gv_i_186;
													for (_gv_i_186 = 0; _gv_i_186 < NUM_OUTPUTS; _gv_i_186 = _gv_i_186 + 1) begin : g_rsp_data_in
														localparam i = _gv_i_186;
														// Trace: src/VX_mem_arb.sv:120:13
														assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_valid;
														// Trace: src/VX_mem_arb.sv:121:13
														assign rsp_data_in[i * 131+:131] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_data;
														// Trace: src/VX_mem_arb.sv:122:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_nc_arb_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
													end
													// Trace: src/VX_mem_arb.sv:124:9
													VX_stream_arb #(
														.NUM_INPUTS(NUM_OUTPUTS),
														.NUM_OUTPUTS(NUM_INPUTS),
														.DATAW(RSP_DATAW),
														.ARBITER(ARBITER),
														.OUT_BUF(RSP_OUT_BUF)
													) req_arb(
														.clk(clk),
														.reset(reset),
														.valid_in(rsp_valid_in),
														.ready_in(rsp_ready_in),
														.data_in(rsp_data_in),
														.data_out(rsp_data_out),
														.valid_out(rsp_valid_out),
														.ready_out(rsp_ready_out),
														.sel_out()
													);
												end
												// Trace: src/VX_mem_arb.sv:142:5
												genvar _gv_i_187;
												for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
													localparam i = _gv_i_187;
													// Trace: src/VX_mem_arb.sv:143:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
													// Trace: src/VX_mem_arb.sv:144:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 131+:131];
													// Trace: src/VX_mem_arb.sv:145:9
													assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.core_bus_in_nc_if[i + _mbase_bus_in_if].rsp_ready;
												end
											end
											assign core_bus_nc_arb.clk = clk;
											assign core_bus_nc_arb.reset = reset;
											// Trace: src/VX_cache_bypass.sv:101:5
											// expanded interface instance: mem_bus_out_nc_if
											localparam _param_0061C_DATA_SIZE = LINE_SIZE;
											localparam _param_0061C_TAG_WIDTH = MEM_TAG_NC2_WIDTH;
											genvar _arr_0061C;
											for (_arr_0061C = 0; _arr_0061C <= 0; _arr_0061C = _arr_0061C + 1) begin : mem_bus_out_nc_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_0061C_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_0061C_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [610:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [516:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache_bypass.sv:105:5
											genvar _gv_i_58;
											localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
											localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
											for (_gv_i_58 = 0; _gv_i_58 < MEM_PORTS; _gv_i_58 = _gv_i_58 + 1) begin : g_mem_bus_out_nc
												localparam i = _gv_i_58;
												// Trace: src/VX_cache_bypass.sv:106:9
												wire core_req_nc_arb_rw;
												// Trace: src/VX_cache_bypass.sv:107:9
												wire [15:0] core_req_nc_arb_byteen;
												// Trace: src/VX_cache_bypass.sv:108:9
												wire [27:0] core_req_nc_arb_addr;
												// Trace: src/VX_cache_bypass.sv:109:9
												wire [2:0] core_req_nc_arb_flags;
												// Trace: src/VX_cache_bypass.sv:110:9
												wire [127:0] core_req_nc_arb_data;
												// Trace: src/VX_cache_bypass.sv:111:9
												wire [2:0] core_req_nc_arb_tag;
												// Trace: src/VX_cache_bypass.sv:112:9
												assign {core_req_nc_arb_rw, core_req_nc_arb_addr, core_req_nc_arb_data, core_req_nc_arb_byteen, core_req_nc_arb_flags, core_req_nc_arb_tag} = core_bus_nc_arb_if[i].req_data;
												// Trace: src/VX_cache_bypass.sv:120:9
												wire [25:0] core_req_nc_arb_addr_w;
												// Trace: src/VX_cache_bypass.sv:121:9
												reg [63:0] core_req_nc_arb_byteen_w;
												// Trace: src/VX_cache_bypass.sv:122:9
												reg [511:0] core_req_nc_arb_data_w;
												// Trace: src/VX_cache_bypass.sv:123:9
												wire [127:0] core_rsp_nc_arb_data_w;
												// Trace: src/VX_cache_bypass.sv:124:9
												wire [4:0] core_req_nc_arb_tag_w;
												// Trace: src/VX_cache_bypass.sv:125:9
												wire [2:0] core_rsp_nc_arb_tag_w;
												if (1) begin : g_multi_word_line
													// Trace: src/VX_cache_bypass.sv:127:13
													wire [1:0] rsp_wsel;
													// Trace: src/VX_cache_bypass.sv:128:13
													wire [1:0] req_wsel = core_req_nc_arb_addr[1:0];
													// Trace: src/VX_cache_bypass.sv:129:13
													always @(*) begin
														// Trace: src/VX_cache_bypass.sv:130:17
														core_req_nc_arb_byteen_w = 1'sb0;
														// Trace: src/VX_cache_bypass.sv:131:17
														core_req_nc_arb_byteen_w[req_wsel * 16+:16] = core_req_nc_arb_byteen;
														// Trace: src/VX_cache_bypass.sv:132:17
														core_req_nc_arb_data_w = 1'sbx;
														// Trace: src/VX_cache_bypass.sv:133:17
														core_req_nc_arb_data_w[req_wsel * 128+:128] = core_req_nc_arb_data;
													end
													// Trace: src/VX_cache_bypass.sv:135:13
													VX_bits_insert #(
														.N(MEM_TAG_NC1_WIDTH),
														.S(WSEL_BITS),
														.POS(TAG_SEL_IDX)
													) wsel_insert(
														.data_in(core_req_nc_arb_tag),
														.ins_in(req_wsel),
														.data_out(core_req_nc_arb_tag_w)
													);
													// Trace: src/VX_cache_bypass.sv:144:13
													VX_bits_remove #(
														.N(MEM_TAG_NC2_WIDTH),
														.S(WSEL_BITS),
														.POS(TAG_SEL_IDX)
													) wsel_remove(
														.data_in(mem_bus_out_nc_if[i].rsp_data[4-:5]),
														.sel_out(rsp_wsel),
														.data_out(core_rsp_nc_arb_tag_w)
													);
													// Trace: src/VX_cache_bypass.sv:153:13
													assign core_req_nc_arb_addr_w = core_req_nc_arb_addr[WSEL_BITS+:MEM_ADDR_WIDTH];
													// Trace: src/VX_cache_bypass.sv:154:13
													assign core_rsp_nc_arb_data_w = mem_bus_out_nc_if[i].rsp_data[5 + (rsp_wsel * CORE_DATA_WIDTH)+:CORE_DATA_WIDTH];
												end
												// Trace: src/VX_cache_bypass.sv:163:9
												assign mem_bus_out_nc_if[i].req_valid = core_bus_nc_arb_if[i].req_valid;
												// Trace: src/VX_cache_bypass.sv:164:9
												assign mem_bus_out_nc_if[i].req_data = {core_req_nc_arb_rw, core_req_nc_arb_addr_w, core_req_nc_arb_data_w, core_req_nc_arb_byteen_w, core_req_nc_arb_flags, core_req_nc_arb_tag_w};
												// Trace: src/VX_cache_bypass.sv:172:9
												assign core_bus_nc_arb_if[i].req_ready = mem_bus_out_nc_if[i].req_ready;
												// Trace: src/VX_cache_bypass.sv:173:9
												assign core_bus_nc_arb_if[i].rsp_valid = mem_bus_out_nc_if[i].rsp_valid;
												// Trace: src/VX_cache_bypass.sv:174:9
												assign core_bus_nc_arb_if[i].rsp_data = {core_rsp_nc_arb_data_w, core_rsp_nc_arb_tag_w};
												// Trace: src/VX_cache_bypass.sv:178:9
												assign mem_bus_out_nc_if[i].rsp_ready = core_bus_nc_arb_if[i].rsp_ready;
											end
											// Trace: src/VX_cache_bypass.sv:180:5
											// expanded interface instance: mem_bus_out_src_if
											localparam _param_913F6_DATA_SIZE = LINE_SIZE;
											localparam _param_913F6_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
											genvar _arr_913F6;
											for (_arr_913F6 = 0; _arr_913F6 <= (((CACHE_ENABLE ? 2 : 1) * MEM_PORTS) - 1); _arr_913F6 = _arr_913F6 + 1) begin : mem_bus_out_src_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_913F6_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_913F6_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [610:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [516:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache_bypass.sv:184:5
											genvar _gv_i_59;
											for (_gv_i_59 = 0; _gv_i_59 < MEM_PORTS; _gv_i_59 = _gv_i_59 + 1) begin : g_mem_bus_out_src
												localparam i = _gv_i_59;
												// Trace: src/VX_cache_bypass.sv:186:5
												assign mem_bus_out_src_if[0 + i].req_valid = mem_bus_out_nc_if[i].req_valid;
												// Trace: src/VX_cache_bypass.sv:187:5
												assign mem_bus_out_src_if[0 + i].req_data[610] = mem_bus_out_nc_if[i].req_data[610];
												// Trace: src/VX_cache_bypass.sv:188:5
												assign mem_bus_out_src_if[0 + i].req_data[609-:26] = mem_bus_out_nc_if[i].req_data[609-:26];
												// Trace: src/VX_cache_bypass.sv:189:5
												assign mem_bus_out_src_if[0 + i].req_data[583-:512] = mem_bus_out_nc_if[i].req_data[583-:512];
												// Trace: src/VX_cache_bypass.sv:190:5
												assign mem_bus_out_src_if[0 + i].req_data[71-:64] = mem_bus_out_nc_if[i].req_data[71-:64];
												// Trace: src/VX_cache_bypass.sv:191:5
												assign mem_bus_out_src_if[0 + i].req_data[7-:3] = mem_bus_out_nc_if[i].req_data[7-:3];
												if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk1
													if (1) begin : genblk1
														if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
															// Trace: src/VX_cache_bypass.sv:195:17
															assign mem_bus_out_src_if[0 + i].req_data[4-:5] = {mem_bus_out_nc_if[i].req_data[4-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_NC2_WIDTH {1'b0}}, mem_bus_out_nc_if[i].req_data[3-:4]};
														end
														else begin : genblk1
															// Trace: src/VX_cache_bypass.sv:197:17
															assign mem_bus_out_src_if[0 + i].req_data[4-:5] = {mem_bus_out_nc_if[i].req_data[4-:1], mem_bus_out_nc_if[i].req_data[(MEM_TAG_OUT_WIDTH - VX_gpu_pkg_UUID_WIDTH) - 1:0]};
														end
													end
												end
												else begin : genblk1
													// Trace: src/VX_cache_bypass.sv:207:9
													assign mem_bus_out_src_if[0 + i].req_data[4-:5] = mem_bus_out_nc_if[i].req_data[4-:5];
												end
												// Trace: src/VX_cache_bypass.sv:209:5
												assign mem_bus_out_nc_if[i].req_ready = mem_bus_out_src_if[0 + i].req_ready;
												// Trace: src/VX_cache_bypass.sv:210:5
												assign mem_bus_out_nc_if[i].rsp_valid = mem_bus_out_src_if[0 + i].rsp_valid;
												// Trace: src/VX_cache_bypass.sv:211:5
												assign mem_bus_out_nc_if[i].rsp_data[516-:512] = mem_bus_out_src_if[0 + i].rsp_data[516-:512];
												if (MEM_TAG_OUT_WIDTH != MEM_TAG_NC2_WIDTH) begin : genblk2
													if (1) begin : genblk1
														if (MEM_TAG_OUT_WIDTH > MEM_TAG_NC2_WIDTH) begin : genblk1
															// Trace: src/VX_cache_bypass.sv:215:17
															assign mem_bus_out_nc_if[i].rsp_data[4-:5] = {mem_bus_out_src_if[0 + i].rsp_data[4-:1], mem_bus_out_src_if[0 + i].rsp_data[3:0]};
														end
														else begin : genblk1
															// Trace: src/VX_cache_bypass.sv:217:17
															assign mem_bus_out_nc_if[i].rsp_data[4-:5] = {mem_bus_out_src_if[0 + i].rsp_data[4-:1], {MEM_TAG_NC2_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[0 + i].rsp_data[3-:4]};
														end
													end
												end
												else begin : genblk2
													// Trace: src/VX_cache_bypass.sv:227:9
													assign mem_bus_out_nc_if[i].rsp_data[4-:5] = mem_bus_out_src_if[0 + i].rsp_data[4-:5];
												end
												// Trace: src/VX_cache_bypass.sv:229:5
												assign mem_bus_out_src_if[0 + i].rsp_ready = mem_bus_out_nc_if[i].rsp_ready;
												if (CACHE_ENABLE) begin : g_cache
													// Trace: src/VX_cache_bypass.sv:233:5
													assign mem_bus_out_src_if[1 + i].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_valid;
													// Trace: src/VX_cache_bypass.sv:234:5
													assign mem_bus_out_src_if[1 + i].req_data[610] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[610];
													// Trace: src/VX_cache_bypass.sv:235:5
													assign mem_bus_out_src_if[1 + i].req_data[609-:26] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[609-:26];
													// Trace: src/VX_cache_bypass.sv:236:5
													assign mem_bus_out_src_if[1 + i].req_data[583-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[583-:512];
													// Trace: src/VX_cache_bypass.sv:237:5
													assign mem_bus_out_src_if[1 + i].req_data[71-:64] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[71-:64];
													// Trace: src/VX_cache_bypass.sv:238:5
													assign mem_bus_out_src_if[1 + i].req_data[7-:3] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[7-:3];
													if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk1
														if (1) begin : genblk1
															if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
																// Trace: src/VX_cache_bypass.sv:242:17
																assign mem_bus_out_src_if[1 + i].req_data[4-:5] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], {MEM_TAG_OUT_WIDTH - MEM_TAG_IN_WIDTH {1'b0}}, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[3-:4]};
															end
															else begin : genblk1
																// Trace: src/VX_cache_bypass.sv:244:17
																assign mem_bus_out_src_if[1 + i].req_data[4-:5] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[(MEM_TAG_OUT_WIDTH - VX_gpu_pkg_UUID_WIDTH) - 1:0]};
															end
														end
													end
													else begin : genblk1
														// Trace: src/VX_cache_bypass.sv:254:9
														assign mem_bus_out_src_if[1 + i].req_data[4-:5] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_data[4-:5];
													end
													// Trace: src/VX_cache_bypass.sv:256:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = mem_bus_out_src_if[1 + i].req_ready;
													// Trace: src/VX_cache_bypass.sv:257:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = mem_bus_out_src_if[1 + i].rsp_valid;
													// Trace: src/VX_cache_bypass.sv:258:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[516-:512] = mem_bus_out_src_if[1 + i].rsp_data[516-:512];
													if (MEM_TAG_OUT_WIDTH != MEM_TAG_IN_WIDTH) begin : genblk2
														if (1) begin : genblk1
															if (MEM_TAG_OUT_WIDTH > MEM_TAG_IN_WIDTH) begin : genblk1
																// Trace: src/VX_cache_bypass.sv:262:17
																assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[4-:1], mem_bus_out_src_if[1 + i].rsp_data[3:0]};
															end
															else begin : genblk1
																// Trace: src/VX_cache_bypass.sv:264:17
																assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = {mem_bus_out_src_if[1 + i].rsp_data[4-:1], {MEM_TAG_IN_WIDTH - MEM_TAG_OUT_WIDTH {1'b0}}, mem_bus_out_src_if[1 + i].rsp_data[3-:4]};
															end
														end
													end
													else begin : genblk2
														// Trace: src/VX_cache_bypass.sv:274:9
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data[4-:5] = mem_bus_out_src_if[1 + i].rsp_data[4-:5];
													end
													// Trace: src/VX_cache_bypass.sv:276:5
													assign mem_bus_out_src_if[1 + i].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_ready;
												end
												else begin : g_no_cache
													// Trace: src/VX_cache_bypass.sv:279:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].req_ready = 0;
													// Trace: src/VX_cache_bypass.sv:280:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_valid = 0;
													// Trace: src/VX_cache_bypass.sv:281:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_in_if].rsp_data = 1'sb0;
												end
											end
											// Trace: src/VX_cache_bypass.sv:284:5
											// expanded module instance: mem_bus_out_arb
											localparam _bbase_B06D0_bus_in_if = 0;
											localparam _bbase_B06D0_bus_out_if = 0;
											localparam _param_B06D0_NUM_INPUTS = (CACHE_ENABLE ? 2 : 1) * MEM_PORTS;
											localparam _param_B06D0_NUM_OUTPUTS = MEM_PORTS;
											localparam _param_B06D0_DATA_SIZE = LINE_SIZE;
											localparam _param_B06D0_TAG_WIDTH = MEM_TAG_OUT_WIDTH;
											localparam _param_B06D0_ARBITER = "R";
											localparam _param_B06D0_REQ_OUT_BUF = (DIRECT_PASSTHRU ? 0 : 2);
											localparam _param_B06D0_RSP_OUT_BUF = 0;
											if (1) begin : mem_bus_out_arb
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_arb.sv:2:15
												localparam NUM_INPUTS = _param_B06D0_NUM_INPUTS;
												// Trace: src/VX_mem_arb.sv:3:15
												localparam NUM_OUTPUTS = _param_B06D0_NUM_OUTPUTS;
												// Trace: src/VX_mem_arb.sv:4:15
												localparam DATA_SIZE = _param_B06D0_DATA_SIZE;
												// Trace: src/VX_mem_arb.sv:5:15
												localparam TAG_WIDTH = _param_B06D0_TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:6:15
												localparam TAG_SEL_IDX = 0;
												// Trace: src/VX_mem_arb.sv:7:15
												localparam REQ_OUT_BUF = _param_B06D0_REQ_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:8:15
												localparam RSP_OUT_BUF = _param_B06D0_RSP_OUT_BUF;
												// Trace: src/VX_mem_arb.sv:9:15
												localparam ARBITER = _param_B06D0_ARBITER;
												// Trace: src/VX_mem_arb.sv:10:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_arb.sv:11:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_arb.sv:12:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_arb.sv:14:5
												wire clk;
												// Trace: src/VX_mem_arb.sv:15:5
												wire reset;
												// Trace: src/VX_mem_arb.sv:16:5
												localparam _mbase_bus_in_if = 0;
												// Trace: src/VX_mem_arb.sv:17:5
												localparam _mbase_bus_out_if = 0;
												// Trace: src/VX_mem_arb.sv:19:5
												localparam DATA_WIDTH = 512;
												// Trace: src/VX_mem_arb.sv:20:5
												localparam LOG_NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? $clog2((NUM_INPUTS + 0) / 1) : 0);
												// Trace: src/VX_mem_arb.sv:21:5
												localparam REQ_DATAW = 606 + TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:22:5
												localparam RSP_DATAW = DATA_WIDTH + TAG_WIDTH;
												// Trace: src/VX_mem_arb.sv:23:5
												localparam SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
												// Trace: src/VX_mem_arb.sv:24:5
												wire [NUM_INPUTS - 1:0] req_valid_in;
												// Trace: src/VX_mem_arb.sv:25:5
												wire [(NUM_INPUTS * REQ_DATAW) - 1:0] req_data_in;
												// Trace: src/VX_mem_arb.sv:26:5
												wire [NUM_INPUTS - 1:0] req_ready_in;
												// Trace: src/VX_mem_arb.sv:27:5
												wire [0:0] req_valid_out;
												// Trace: src/VX_mem_arb.sv:28:5
												wire [REQ_DATAW - 1:0] req_data_out;
												// Trace: src/VX_mem_arb.sv:29:5
												wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] req_sel_out;
												// Trace: src/VX_mem_arb.sv:30:5
												wire [0:0] req_ready_out;
												// Trace: src/VX_mem_arb.sv:31:5
												genvar _gv_i_183;
												for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
													localparam i = _gv_i_183;
													// Trace: src/VX_mem_arb.sv:32:9
													assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_valid;
													// Trace: src/VX_mem_arb.sv:33:9
													assign req_data_in[i * 611+:611] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_data;
													// Trace: src/VX_mem_arb.sv:34:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
												end
												// Trace: src/VX_mem_arb.sv:36:5
												VX_stream_arb #(
													.NUM_INPUTS(NUM_INPUTS),
													.NUM_OUTPUTS(NUM_OUTPUTS),
													.DATAW(REQ_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(REQ_OUT_BUF)
												) req_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(req_valid_in),
													.ready_in(req_ready_in),
													.data_in(req_data_in),
													.data_out(req_data_out),
													.sel_out(req_sel_out),
													.valid_out(req_valid_out),
													.ready_out(req_ready_out)
												);
												// Trace: src/VX_mem_arb.sv:53:5
												genvar _gv_i_184;
												for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
													localparam i = _gv_i_184;
													// Trace: src/VX_mem_arb.sv:54:9
													wire [TAG_WIDTH - 1:0] req_tag_out;
													// Trace: src/VX_mem_arb.sv:55:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
													// Trace: src/VX_mem_arb.sv:56:9
													assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[611], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[610-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[584-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[72-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[8-:3], req_tag_out} = req_data_out[i * 611+:611];
													// Trace: src/VX_mem_arb.sv:64:9
													assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
													if (NUM_INPUTS > NUM_OUTPUTS) begin : g_req_tag_sel_out
														// Trace: src/VX_mem_arb.sv:66:13
														VX_bits_insert #(
															.N(TAG_WIDTH),
															.S(LOG_NUM_REQS),
															.POS(TAG_SEL_IDX)
														) bits_insert(
															.data_in(req_tag_out),
															.ins_in(req_sel_out[i * 1+:1]),
															.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[5-:6])
														);
													end
													else begin : g_req_tag_out
														// Trace: src/VX_mem_arb.sv:76:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[5-:6] = req_tag_out;
													end
												end
												// Trace: src/VX_mem_arb.sv:79:5
												wire [NUM_INPUTS - 1:0] rsp_valid_out;
												// Trace: src/VX_mem_arb.sv:80:5
												wire [(NUM_INPUTS * RSP_DATAW) - 1:0] rsp_data_out;
												// Trace: src/VX_mem_arb.sv:81:5
												wire [NUM_INPUTS - 1:0] rsp_ready_out;
												// Trace: src/VX_mem_arb.sv:82:5
												wire [0:0] rsp_valid_in;
												// Trace: src/VX_mem_arb.sv:83:5
												wire [RSP_DATAW - 1:0] rsp_data_in;
												// Trace: src/VX_mem_arb.sv:84:5
												wire [0:0] rsp_ready_in;
												// Trace: src/VX_mem_arb.sv:85:5
												if (NUM_INPUTS > NUM_OUTPUTS) begin : g_rsp_select
													// Trace: src/VX_mem_arb.sv:86:9
													wire [LOG_NUM_REQS - 1:0] rsp_sel_in;
													genvar _gv_i_185;
													for (_gv_i_185 = 0; _gv_i_185 < NUM_OUTPUTS; _gv_i_185 = _gv_i_185 + 1) begin : g_rsp_data_in
														localparam i = _gv_i_185;
														// Trace: src/VX_mem_arb.sv:88:13
														wire [TAG_WIDTH - 1:0] rsp_tag_out;
														// Trace: src/VX_mem_arb.sv:89:13
														VX_bits_remove #(
															.N(TAG_WIDTH + LOG_NUM_REQS),
															.S(LOG_NUM_REQS),
															.POS(TAG_SEL_IDX)
														) bits_remove(
															.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[5-:6]),
															.sel_out(rsp_sel_in[i * 1+:1]),
															.data_out(rsp_tag_out)
														);
														// Trace: src/VX_mem_arb.sv:98:13
														assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
														// Trace: src/VX_mem_arb.sv:99:13
														assign rsp_data_in[i * 517+:517] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data[517-:512], rsp_tag_out};
														// Trace: src/VX_mem_arb.sv:100:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
													end
													// Trace: src/VX_mem_arb.sv:102:9
													VX_stream_switch #(
														.NUM_INPUTS(NUM_OUTPUTS),
														.NUM_OUTPUTS(NUM_INPUTS),
														.DATAW(RSP_DATAW),
														.OUT_BUF(RSP_OUT_BUF)
													) rsp_switch(
														.clk(clk),
														.reset(reset),
														.sel_in(rsp_sel_in),
														.valid_in(rsp_valid_in),
														.ready_in(rsp_ready_in),
														.data_in(rsp_data_in),
														.data_out(rsp_data_out),
														.valid_out(rsp_valid_out),
														.ready_out(rsp_ready_out)
													);
												end
												else begin : g_rsp_arb
													genvar _gv_i_186;
													for (_gv_i_186 = 0; _gv_i_186 < NUM_OUTPUTS; _gv_i_186 = _gv_i_186 + 1) begin : g_rsp_data_in
														localparam i = _gv_i_186;
														// Trace: src/VX_mem_arb.sv:120:13
														assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
														// Trace: src/VX_mem_arb.sv:121:13
														assign rsp_data_in[i * 517+:517] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
														// Trace: src/VX_mem_arb.sv:122:13
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
													end
													// Trace: src/VX_mem_arb.sv:124:9
													VX_stream_arb #(
														.NUM_INPUTS(NUM_OUTPUTS),
														.NUM_OUTPUTS(NUM_INPUTS),
														.DATAW(RSP_DATAW),
														.ARBITER(ARBITER),
														.OUT_BUF(RSP_OUT_BUF)
													) req_arb(
														.clk(clk),
														.reset(reset),
														.valid_in(rsp_valid_in),
														.ready_in(rsp_ready_in),
														.data_in(rsp_data_in),
														.data_out(rsp_data_out),
														.valid_out(rsp_valid_out),
														.ready_out(rsp_ready_out),
														.sel_out()
													);
												end
												// Trace: src/VX_mem_arb.sv:142:5
												genvar _gv_i_187;
												for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
													localparam i = _gv_i_187;
													// Trace: src/VX_mem_arb.sv:143:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
													// Trace: src/VX_mem_arb.sv:144:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 517+:517];
													// Trace: src/VX_mem_arb.sv:145:9
													assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_bypass.cache_bypass.mem_bus_out_src_if[i + _mbase_bus_in_if].rsp_ready;
												end
											end
											assign mem_bus_out_arb.clk = clk;
											assign mem_bus_out_arb.reset = reset;
										end
										assign cache_bypass.clk = clk;
										assign cache_bypass.reset = reset;
									end
									else begin : g_no_bypass
										genvar _gv_i_38;
										for (_gv_i_38 = 0; _gv_i_38 < NUM_REQS; _gv_i_38 = _gv_i_38 + 1) begin : g_core_bus_cache_if
											localparam i = _gv_i_38;
											// Trace: src/VX_cache_wrap.sv:73:5
											assign core_bus_cache_if[i].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_if].req_valid;
											// Trace: src/VX_cache_wrap.sv:74:5
											assign core_bus_cache_if[i].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_if].req_data;
											// Trace: src/VX_cache_wrap.sv:75:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_if].req_ready = core_bus_cache_if[i].req_ready;
											// Trace: src/VX_cache_wrap.sv:76:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_if].rsp_valid = core_bus_cache_if[i].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:77:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_if].rsp_data = core_bus_cache_if[i].rsp_data;
											// Trace: src/VX_cache_wrap.sv:78:5
											assign core_bus_cache_if[i].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.arb_core_bus_if[i + _mbase_core_bus_if].rsp_ready;
										end
										genvar _gv_i_39;
										for (_gv_i_39 = 0; _gv_i_39 < MEM_PORTS; _gv_i_39 = _gv_i_39 + 1) begin : g_mem_bus_tmp_if
											localparam i = _gv_i_39;
											// Trace: src/VX_cache_wrap.sv:81:5
											assign mem_bus_tmp_if[i].req_valid = mem_bus_cache_if[i].req_valid;
											// Trace: src/VX_cache_wrap.sv:82:5
											assign mem_bus_tmp_if[i].req_data = mem_bus_cache_if[i].req_data;
											// Trace: src/VX_cache_wrap.sv:83:5
											assign mem_bus_cache_if[i].req_ready = mem_bus_tmp_if[i].req_ready;
											// Trace: src/VX_cache_wrap.sv:84:5
											assign mem_bus_cache_if[i].rsp_valid = mem_bus_tmp_if[i].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:85:5
											assign mem_bus_cache_if[i].rsp_data = mem_bus_tmp_if[i].rsp_data;
											// Trace: src/VX_cache_wrap.sv:86:5
											assign mem_bus_tmp_if[i].rsp_ready = mem_bus_cache_if[i].rsp_ready;
										end
									end
									// Trace: src/VX_cache_wrap.sv:89:5
									genvar _gv_i_40;
									for (_gv_i_40 = 0; _gv_i_40 < MEM_PORTS; _gv_i_40 = _gv_i_40 + 1) begin : g_mem_bus_if
										localparam i = _gv_i_40;
										if (WRITE_ENABLE) begin : g_we
											// Trace: src/VX_cache_wrap.sv:91:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
											// Trace: src/VX_cache_wrap.sv:92:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[i].req_data;
											// Trace: src/VX_cache_wrap.sv:93:5
											assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
											// Trace: src/VX_cache_wrap.sv:94:5
											assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:95:5
											assign mem_bus_tmp_if[i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
											// Trace: src/VX_cache_wrap.sv:96:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
										end
										else begin : g_ro
											// Trace: src/VX_cache_wrap.sv:98:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
											// Trace: src/VX_cache_wrap.sv:99:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[611] = 0;
											// Trace: src/VX_cache_wrap.sv:100:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[610-:26] = mem_bus_tmp_if[i].req_data[610-:26];
											// Trace: src/VX_cache_wrap.sv:101:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[584-:512] = 1'sb0;
											// Trace: src/VX_cache_wrap.sv:102:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[72-:64] = 1'sb1;
											// Trace: src/VX_cache_wrap.sv:103:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[8-:3] = mem_bus_tmp_if[i].req_data[8-:3];
											// Trace: src/VX_cache_wrap.sv:104:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_data[5-:6] = mem_bus_tmp_if[i].req_data[5-:6];
											// Trace: src/VX_cache_wrap.sv:105:5
											assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
											// Trace: src/VX_cache_wrap.sv:106:5
											assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
											// Trace: src/VX_cache_wrap.sv:107:5
											assign mem_bus_tmp_if[i].rsp_data[517-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[517-:512];
											// Trace: src/VX_cache_wrap.sv:108:5
											assign mem_bus_tmp_if[i].rsp_data[5-:6] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[5-:6];
											// Trace: src/VX_cache_wrap.sv:109:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.cache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
										end
									end
									// Trace: src/VX_cache_wrap.sv:112:5
									if (1) begin : g_cache
										// Trace: src/VX_cache_wrap.sv:113:9
										// expanded module instance: cache
										localparam _bbase_90EE2_core_bus_if = 0;
										localparam _bbase_90EE2_mem_bus_if = 0;
										localparam _param_90EE2_INSTANCE_ID = INSTANCE_ID;
										localparam _param_90EE2_CACHE_SIZE = CACHE_SIZE;
										localparam _param_90EE2_LINE_SIZE = LINE_SIZE;
										localparam _param_90EE2_NUM_BANKS = NUM_BANKS;
										localparam _param_90EE2_NUM_WAYS = NUM_WAYS;
										localparam _param_90EE2_WORD_SIZE = WORD_SIZE;
										localparam _param_90EE2_NUM_REQS = NUM_REQS;
										localparam _param_90EE2_MEM_PORTS = MEM_PORTS;
										localparam _param_90EE2_WRITE_ENABLE = WRITE_ENABLE;
										localparam _param_90EE2_WRITEBACK = WRITEBACK;
										localparam _param_90EE2_DIRTY_BYTES = DIRTY_BYTES;
										localparam _param_90EE2_REPL_POLICY = REPL_POLICY;
										localparam _param_90EE2_CRSQ_SIZE = CRSQ_SIZE;
										localparam _param_90EE2_MSHR_SIZE = MSHR_SIZE;
										localparam _param_90EE2_MRSQ_SIZE = MRSQ_SIZE;
										localparam _param_90EE2_MREQ_SIZE = MREQ_SIZE;
										localparam _param_90EE2_TAG_WIDTH = TAG_WIDTH;
										localparam _param_90EE2_CORE_OUT_BUF = (BYPASS_ENABLE ? 1 : CORE_OUT_BUF);
										localparam _param_90EE2_MEM_OUT_BUF = (BYPASS_ENABLE ? 1 : MEM_OUT_BUF);
										if (1) begin : cache
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_cache.sv:2:15
											localparam INSTANCE_ID = _param_90EE2_INSTANCE_ID;
											// Trace: src/VX_cache.sv:3:15
											localparam NUM_REQS = _param_90EE2_NUM_REQS;
											// Trace: src/VX_cache.sv:4:15
											localparam MEM_PORTS = _param_90EE2_MEM_PORTS;
											// Trace: src/VX_cache.sv:5:15
											localparam CACHE_SIZE = _param_90EE2_CACHE_SIZE;
											// Trace: src/VX_cache.sv:6:15
											localparam LINE_SIZE = _param_90EE2_LINE_SIZE;
											// Trace: src/VX_cache.sv:7:15
											localparam NUM_BANKS = _param_90EE2_NUM_BANKS;
											// Trace: src/VX_cache.sv:8:15
											localparam NUM_WAYS = _param_90EE2_NUM_WAYS;
											// Trace: src/VX_cache.sv:9:15
											localparam WORD_SIZE = _param_90EE2_WORD_SIZE;
											// Trace: src/VX_cache.sv:10:15
											localparam CRSQ_SIZE = _param_90EE2_CRSQ_SIZE;
											// Trace: src/VX_cache.sv:11:15
											localparam MSHR_SIZE = _param_90EE2_MSHR_SIZE;
											// Trace: src/VX_cache.sv:12:15
											localparam MRSQ_SIZE = _param_90EE2_MRSQ_SIZE;
											// Trace: src/VX_cache.sv:13:15
											localparam MREQ_SIZE = _param_90EE2_MREQ_SIZE;
											// Trace: src/VX_cache.sv:14:15
											localparam WRITE_ENABLE = _param_90EE2_WRITE_ENABLE;
											// Trace: src/VX_cache.sv:15:15
											localparam WRITEBACK = _param_90EE2_WRITEBACK;
											// Trace: src/VX_cache.sv:16:15
											localparam DIRTY_BYTES = _param_90EE2_DIRTY_BYTES;
											// Trace: src/VX_cache.sv:17:15
											localparam REPL_POLICY = _param_90EE2_REPL_POLICY;
											// Trace: src/VX_cache.sv:18:15
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam TAG_WIDTH = _param_90EE2_TAG_WIDTH;
											// Trace: src/VX_cache.sv:19:15
											localparam CORE_OUT_BUF = _param_90EE2_CORE_OUT_BUF;
											// Trace: src/VX_cache.sv:20:15
											localparam MEM_OUT_BUF = _param_90EE2_MEM_OUT_BUF;
											// Trace: src/VX_cache.sv:22:5
											wire clk;
											// Trace: src/VX_cache.sv:23:5
											wire reset;
											// Trace: src/VX_cache.sv:24:5
											localparam _mbase_core_bus_if = 0;
											// Trace: src/VX_cache.sv:25:5
											localparam _mbase_mem_bus_if = 0;
											// Trace: src/VX_cache.sv:27:5
											localparam REQ_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:28:5
											localparam WORD_SEL_WIDTH = 2;
											// Trace: src/VX_cache.sv:29:5
											localparam MSHR_ADDR_WIDTH = 4;
											// Trace: src/VX_cache.sv:30:5
											localparam MEM_TAG_WIDTH = 5;
											// Trace: src/VX_cache.sv:32:5
											localparam WORDS_PER_LINE = 4;
											// Trace: src/VX_cache.sv:33:5
											localparam WORD_WIDTH = 128;
											// Trace: src/VX_cache.sv:34:5
											localparam WORD_SEL_BITS = 2;
											// Trace: src/VX_cache.sv:35:5
											localparam BANK_SEL_BITS = 0;
											// Trace: src/VX_cache.sv:36:5
											localparam BANK_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:37:5
											localparam LINE_ADDR_WIDTH = 26;
											// Trace: src/VX_cache.sv:38:5
											localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
											localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
											localparam CORE_REQ_DATAW = 179;
											// Trace: src/VX_cache.sv:39:5
											localparam CORE_RSP_DATAW = 131;
											// Trace: src/VX_cache.sv:40:5
											localparam BANK_MEM_TAG_WIDTH = 5;
											// Trace: src/VX_cache.sv:41:5
											localparam MEM_REQ_DATAW = 611;
											// Trace: src/VX_cache.sv:42:5
											localparam MEM_RSP_DATAW = 517;
											// Trace: src/VX_cache.sv:43:5
											localparam MEM_PORTS_SEL_BITS = 0;
											// Trace: src/VX_cache.sv:44:5
											localparam MEM_PORTS_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:45:5
											localparam MEM_ARB_SEL_BITS = 0;
											// Trace: src/VX_cache.sv:46:5
											localparam MEM_ARB_SEL_WIDTH = 1;
											// Trace: src/VX_cache.sv:47:5
											localparam REQ_XBAR_BUF = 0;
											// Trace: src/VX_cache.sv:48:5
											localparam CORE_RSP_BUF_ENABLE = 1'd0;
											// Trace: src/VX_cache.sv:49:5
											localparam MEM_REQ_BUF_ENABLE = 1'd0;
											// Trace: src/VX_cache.sv:50:5
											// expanded interface instance: core_bus2_if
											localparam _param_9260A_DATA_SIZE = WORD_SIZE;
											localparam _param_9260A_TAG_WIDTH = TAG_WIDTH;
											genvar _arr_9260A;
											for (_arr_9260A = 0; _arr_9260A <= 0; _arr_9260A = _arr_9260A + 1) begin : core_bus2_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_9260A_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_9260A_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 28;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [178:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [130:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache.sv:54:5
											wire [0:0] per_bank_flush_begin;
											// Trace: src/VX_cache.sv:55:5
											wire [0:0] flush_uuid;
											// Trace: src/VX_cache.sv:56:5
											wire [0:0] per_bank_flush_end;
											// Trace: src/VX_cache.sv:57:5
											wire [0:0] per_bank_core_req_fire;
											// Trace: src/VX_cache.sv:58:5
											// expanded module instance: cache_init
											localparam _bbase_3B3F2_core_bus_in_if = 0;
											localparam _bbase_3B3F2_core_bus_out_if = 0;
											localparam _param_3B3F2_NUM_REQS = NUM_REQS;
											localparam _param_3B3F2_NUM_BANKS = NUM_BANKS;
											localparam _param_3B3F2_TAG_WIDTH = TAG_WIDTH;
											localparam _param_3B3F2_BANK_SEL_LATENCY = 0;
											if (1) begin : cache_init
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_cache_init.sv:2:15
												localparam NUM_REQS = _param_3B3F2_NUM_REQS;
												// Trace: src/VX_cache_init.sv:3:15
												localparam NUM_BANKS = _param_3B3F2_NUM_BANKS;
												// Trace: src/VX_cache_init.sv:4:15
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam TAG_WIDTH = _param_3B3F2_TAG_WIDTH;
												// Trace: src/VX_cache_init.sv:5:15
												localparam BANK_SEL_LATENCY = _param_3B3F2_BANK_SEL_LATENCY;
												// Trace: src/VX_cache_init.sv:7:5
												wire clk;
												// Trace: src/VX_cache_init.sv:8:5
												wire reset;
												// Trace: src/VX_cache_init.sv:9:5
												localparam _mbase_core_bus_in_if = 0;
												// Trace: src/VX_cache_init.sv:10:5
												localparam _mbase_core_bus_out_if = 0;
												// Trace: src/VX_cache_init.sv:11:5
												wire [0:0] bank_req_fire;
												// Trace: src/VX_cache_init.sv:12:5
												wire [0:0] flush_begin;
												// Trace: src/VX_cache_init.sv:13:5
												wire [0:0] flush_uuid;
												// Trace: src/VX_cache_init.sv:14:5
												wire [0:0] flush_end;
												// Trace: src/VX_cache_init.sv:16:5
												localparam STATE_IDLE = 0;
												// Trace: src/VX_cache_init.sv:17:5
												localparam STATE_WAIT1 = 1;
												// Trace: src/VX_cache_init.sv:18:5
												localparam STATE_FLUSH = 2;
												// Trace: src/VX_cache_init.sv:19:5
												localparam STATE_WAIT2 = 3;
												// Trace: src/VX_cache_init.sv:20:5
												localparam STATE_DONE = 4;
												// Trace: src/VX_cache_init.sv:21:5
												reg [2:0] state;
												reg [2:0] state_n;
												// Trace: src/VX_cache_init.sv:22:5
												wire no_inflight_reqs;
												// Trace: src/VX_cache_init.sv:23:5
												if (1) begin : g_no_bank_sel_latency
													// Trace: src/VX_cache_init.sv:62:9
													assign no_inflight_reqs = 0;
												end
												// Trace: src/VX_cache_init.sv:64:5
												reg [0:0] flush_done;
												reg [0:0] flush_done_n;
												// Trace: src/VX_cache_init.sv:65:5
												wire [0:0] flush_req_mask;
												// Trace: src/VX_cache_init.sv:66:5
												genvar _gv_i_215;
												localparam VX_gpu_pkg_MEM_REQ_FLAG_FLUSH = 0;
												for (_gv_i_215 = 0; _gv_i_215 < NUM_REQS; _gv_i_215 = _gv_i_215 + 1) begin : g_flush_req_mask
													localparam i = _gv_i_215;
													// Trace: src/VX_cache_init.sv:67:9
													assign flush_req_mask[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_data[3];
												end
												// Trace: src/VX_cache_init.sv:69:5
												wire flush_req_enable = |flush_req_mask;
												// Trace: src/VX_cache_init.sv:70:5
												reg [0:0] lock_released;
												reg [0:0] lock_released_n;
												// Trace: src/VX_cache_init.sv:71:5
												reg [0:0] flush_uuid_r;
												reg [0:0] flush_uuid_n;
												// Trace: src/VX_cache_init.sv:72:5
												genvar _gv_i_216;
												for (_gv_i_216 = 0; _gv_i_216 < NUM_REQS; _gv_i_216 = _gv_i_216 + 1) begin : g_core_bus_out_req
													localparam i = _gv_i_216;
													// Trace: src/VX_cache_init.sv:73:9
													wire input_enable = ~flush_req_enable || lock_released[i];
													// Trace: src/VX_cache_init.sv:74:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_valid && input_enable;
													// Trace: src/VX_cache_init.sv:75:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_data;
													// Trace: src/VX_cache_init.sv:76:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_ready && input_enable;
												end
												// Trace: src/VX_cache_init.sv:78:5
												genvar _gv_i_217;
												for (_gv_i_217 = 0; _gv_i_217 < NUM_REQS; _gv_i_217 = _gv_i_217 + 1) begin : g_core_bus_in_rsp
													localparam i = _gv_i_217;
													// Trace: src/VX_cache_init.sv:79:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].rsp_valid;
													// Trace: src/VX_cache_init.sv:80:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].rsp_data;
													// Trace: src/VX_cache_init.sv:81:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].rsp_ready;
												end
												// Trace: src/VX_cache_init.sv:83:5
												reg [0:0] core_bus_out_uuid;
												// Trace: src/VX_cache_init.sv:84:5
												wire [0:0] core_bus_out_ready;
												// Trace: src/VX_cache_init.sv:85:5
												genvar _gv_i_218;
												for (_gv_i_218 = 0; _gv_i_218 < NUM_REQS; _gv_i_218 = _gv_i_218 + 1) begin : g_core_bus_out_uuid
													localparam i = _gv_i_218;
													if (1) begin : g_uuid
														// Trace: src/VX_cache_init.sv:87:13
														wire [1:1] sv2v_tmp_FD406;
														assign sv2v_tmp_FD406 = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.core_bus_cache_if[i + _mbase_core_bus_in_if].req_data[2-:1];
														always @(*) core_bus_out_uuid[i+:1] = sv2v_tmp_FD406;
													end
												end
												// Trace: src/VX_cache_init.sv:92:5
												genvar _gv_i_219;
												for (_gv_i_219 = 0; _gv_i_219 < NUM_REQS; _gv_i_219 = _gv_i_219 + 1) begin : g_core_bus_out_ready
													localparam i = _gv_i_219;
													// Trace: src/VX_cache_init.sv:93:9
													assign core_bus_out_ready[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.g_cache.cache.core_bus2_if[i + _mbase_core_bus_out_if].req_ready;
												end
												// Trace: src/VX_cache_init.sv:95:5
												always @(*) begin
													// Trace: src/VX_cache_init.sv:96:9
													state_n = state;
													// Trace: src/VX_cache_init.sv:97:9
													flush_done_n = flush_done;
													// Trace: src/VX_cache_init.sv:98:9
													lock_released_n = lock_released;
													// Trace: src/VX_cache_init.sv:99:9
													flush_uuid_n = flush_uuid_r;
													// Trace: src/VX_cache_init.sv:100:9
													case (state)
														default:
															// Trace: src/VX_cache_init.sv:102:17
															if (flush_req_enable) begin
																// Trace: src/VX_cache_init.sv:103:21
																state_n = STATE_FLUSH;
																// Trace: src/VX_cache_init.sv:104:21
																begin : sv2v_autoblock_2
																	// Trace: src/VX_cache_init.sv:104:26
																	integer i;
																	// Trace: src/VX_cache_init.sv:104:26
																	for (i = 0; i >= 0; i = i - 1)
																		begin
																			// Trace: src/VX_cache_init.sv:105:25
																			if (flush_req_mask[i])
																				// Trace: src/VX_cache_init.sv:106:29
																				flush_uuid_n = core_bus_out_uuid[i+:1];
																		end
																end
															end
														STATE_WAIT1:
															// Trace: src/VX_cache_init.sv:112:17
															if (no_inflight_reqs)
																// Trace: src/VX_cache_init.sv:113:21
																state_n = STATE_FLUSH;
														STATE_FLUSH:
															// Trace: src/VX_cache_init.sv:117:17
															state_n = STATE_WAIT2;
														STATE_WAIT2: begin
															// Trace: src/VX_cache_init.sv:120:17
															flush_done_n = flush_done | flush_end;
															// Trace: src/VX_cache_init.sv:121:17
															if (flush_done_n == {NUM_BANKS {1'b1}}) begin
																// Trace: src/VX_cache_init.sv:122:21
																state_n = STATE_DONE;
																// Trace: src/VX_cache_init.sv:123:21
																flush_done_n = 1'sb0;
																// Trace: src/VX_cache_init.sv:124:21
																lock_released_n = flush_req_mask;
															end
														end
														STATE_DONE: begin
															// Trace: src/VX_cache_init.sv:128:17
															lock_released_n = lock_released & ~core_bus_out_ready;
															// Trace: src/VX_cache_init.sv:129:17
															if (lock_released_n == 0)
																// Trace: src/VX_cache_init.sv:130:21
																state_n = STATE_IDLE;
														end
													endcase
												end
												// Trace: src/VX_cache_init.sv:135:5
												always @(posedge clk) begin
													// Trace: src/VX_cache_init.sv:136:9
													if (reset) begin
														// Trace: src/VX_cache_init.sv:137:13
														state <= STATE_IDLE;
														// Trace: src/VX_cache_init.sv:138:13
														flush_done <= 1'sb0;
														// Trace: src/VX_cache_init.sv:139:13
														lock_released <= 1'sb0;
													end
													else begin
														// Trace: src/VX_cache_init.sv:141:13
														state <= state_n;
														// Trace: src/VX_cache_init.sv:142:13
														flush_done <= flush_done_n;
														// Trace: src/VX_cache_init.sv:143:13
														lock_released <= lock_released_n;
													end
													// Trace: src/VX_cache_init.sv:145:9
													flush_uuid_r <= flush_uuid_n;
												end
												// Trace: src/VX_cache_init.sv:147:5
												assign flush_begin = {NUM_BANKS {state == STATE_FLUSH}};
												// Trace: src/VX_cache_init.sv:148:5
												assign flush_uuid = flush_uuid_r;
											end
											assign cache_init.clk = clk;
											assign cache_init.reset = reset;
											assign cache_init.bank_req_fire = per_bank_core_req_fire;
											assign per_bank_flush_begin = cache_init.flush_begin;
											assign flush_uuid = cache_init.flush_uuid;
											assign cache_init.flush_end = per_bank_flush_end;
											// Trace: src/VX_cache.sv:73:5
											// expanded interface instance: mem_bus_tmp_if
											localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
											localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH;
											genvar _arr_4FE36;
											for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_mem_bus_if.sv:2:15
												localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
												// Trace: src/VX_mem_bus_if.sv:3:15
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:4:15
												localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
												// Trace: src/VX_mem_bus_if.sv:5:15
												localparam MEM_ADDR_WIDTH = 32;
												// Trace: src/VX_mem_bus_if.sv:6:15
												localparam ADDR_WIDTH = 26;
												// Trace: src/VX_mem_bus_if.sv:8:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type tag_t
												// Trace: src/VX_mem_bus_if.sv:12:5
												// removed localparam type req_data_t
												// Trace: src/VX_mem_bus_if.sv:20:5
												// removed localparam type rsp_data_t
												// Trace: src/VX_mem_bus_if.sv:24:5
												wire req_valid;
												// Trace: src/VX_mem_bus_if.sv:25:5
												wire [610:0] req_data;
												// Trace: src/VX_mem_bus_if.sv:26:5
												wire req_ready;
												// Trace: src/VX_mem_bus_if.sv:27:5
												wire rsp_valid;
												// Trace: src/VX_mem_bus_if.sv:28:5
												wire [516:0] rsp_data;
												// Trace: src/VX_mem_bus_if.sv:29:5
												wire rsp_ready;
												// Trace: src/VX_mem_bus_if.sv:30:5
												// Trace: src/VX_mem_bus_if.sv:38:5
											end
											// Trace: src/VX_cache.sv:77:5
											wire [0:0] mem_rsp_queue_valid;
											// Trace: src/VX_cache.sv:78:5
											wire [516:0] mem_rsp_queue_data;
											// Trace: src/VX_cache.sv:79:5
											wire [0:0] mem_rsp_queue_ready;
											// Trace: src/VX_cache.sv:80:5
											genvar _gv_i_228;
											for (_gv_i_228 = 0; _gv_i_228 < MEM_PORTS; _gv_i_228 = _gv_i_228 + 1) begin : g_mem_rsp_queue
												localparam i = _gv_i_228;
												// Trace: src/VX_cache.sv:81:9
												VX_elastic_buffer #(
													.DATAW(MEM_RSP_DATAW),
													.SIZE(MRSQ_SIZE),
													.OUT_REG(1'd1)
												) mem_rsp_queue(
													.clk(clk),
													.reset(reset),
													.valid_in(mem_bus_tmp_if[i].rsp_valid),
													.data_in(mem_bus_tmp_if[i].rsp_data),
													.ready_in(mem_bus_tmp_if[i].rsp_ready),
													.valid_out(mem_rsp_queue_valid[i]),
													.data_out(mem_rsp_queue_data[i * 517+:517]),
													.ready_out(mem_rsp_queue_ready[i])
												);
											end
											// Trace: src/VX_cache.sv:96:5
											wire [516:0] mem_rsp_queue_data_s;
											// Trace: src/VX_cache.sv:97:5
											wire [0:0] mem_rsp_queue_sel;
											// Trace: src/VX_cache.sv:98:5
											genvar _gv_i_229;
											for (_gv_i_229 = 0; _gv_i_229 < MEM_PORTS; _gv_i_229 = _gv_i_229 + 1) begin : g_mem_rsp_queue_data_s
												localparam i = _gv_i_229;
												// Trace: src/VX_cache.sv:99:9
												wire [4:0] mem_rsp_tag_s = mem_rsp_queue_data[(i * 517) + 4-:5];
												// Trace: src/VX_cache.sv:100:9
												wire [511:0] mem_rsp_data_s = mem_rsp_queue_data[(i * 517) + 516-:512];
												// Trace: src/VX_cache.sv:101:9
												assign mem_rsp_queue_data_s[i * 517+:517] = {mem_rsp_data_s, mem_rsp_tag_s};
											end
											// Trace: src/VX_cache.sv:103:5
											genvar _gv_i_230;
											for (_gv_i_230 = 0; _gv_i_230 < MEM_PORTS; _gv_i_230 = _gv_i_230 + 1) begin : g_mem_rsp_queue_sel
												localparam i = _gv_i_230;
												if (1) begin : g_singlebank
													// Trace: src/VX_cache.sv:118:13
													assign mem_rsp_queue_sel[i+:1] = 0;
												end
											end
											// Trace: src/VX_cache.sv:121:5
											wire [0:0] per_bank_mem_rsp_valid;
											// Trace: src/VX_cache.sv:122:5
											wire [516:0] per_bank_mem_rsp_pdata;
											// Trace: src/VX_cache.sv:123:5
											wire [0:0] per_bank_mem_rsp_ready;
											// Trace: src/VX_cache.sv:124:5
											VX_stream_omega #(
												.NUM_INPUTS(MEM_PORTS),
												.NUM_OUTPUTS(NUM_BANKS),
												.DATAW(517),
												.ARBITER("R"),
												.OUT_BUF(3)
											) mem_rsp_xbar(
												.clk(clk),
												.reset(reset),
												.valid_in(mem_rsp_queue_valid),
												.data_in(mem_rsp_queue_data_s),
												.sel_in(mem_rsp_queue_sel),
												.ready_in(mem_rsp_queue_ready),
												.valid_out(per_bank_mem_rsp_valid),
												.data_out(per_bank_mem_rsp_pdata),
												.sel_out(),
												.ready_out(per_bank_mem_rsp_ready),
												.collisions()
											);
											// Trace: src/VX_cache.sv:143:5
											wire [511:0] per_bank_mem_rsp_data;
											// Trace: src/VX_cache.sv:144:5
											wire [4:0] per_bank_mem_rsp_tag;
											// Trace: src/VX_cache.sv:145:5
											genvar _gv_i_231;
											for (_gv_i_231 = 0; _gv_i_231 < NUM_BANKS; _gv_i_231 = _gv_i_231 + 1) begin : g_per_bank_mem_rsp_data
												localparam i = _gv_i_231;
												// Trace: src/VX_cache.sv:146:9
												assign {per_bank_mem_rsp_data[i * 512+:512], per_bank_mem_rsp_tag[i * 5+:5]} = per_bank_mem_rsp_pdata[i * 517+:517];
											end
											// Trace: src/VX_cache.sv:151:5
											wire [0:0] per_bank_core_req_valid;
											// Trace: src/VX_cache.sv:152:5
											wire [25:0] per_bank_core_req_addr;
											// Trace: src/VX_cache.sv:153:5
											wire [0:0] per_bank_core_req_rw;
											// Trace: src/VX_cache.sv:154:5
											wire [1:0] per_bank_core_req_wsel;
											// Trace: src/VX_cache.sv:155:5
											wire [15:0] per_bank_core_req_byteen;
											// Trace: src/VX_cache.sv:156:5
											wire [127:0] per_bank_core_req_data;
											// Trace: src/VX_cache.sv:157:5
											wire [2:0] per_bank_core_req_tag;
											// Trace: src/VX_cache.sv:158:5
											wire [0:0] per_bank_core_req_idx;
											// Trace: src/VX_cache.sv:159:5
											wire [2:0] per_bank_core_req_flags;
											// Trace: src/VX_cache.sv:160:5
											wire [0:0] per_bank_core_req_ready;
											// Trace: src/VX_cache.sv:161:5
											wire [0:0] per_bank_core_rsp_valid;
											// Trace: src/VX_cache.sv:162:5
											wire [127:0] per_bank_core_rsp_data;
											// Trace: src/VX_cache.sv:163:5
											wire [2:0] per_bank_core_rsp_tag;
											// Trace: src/VX_cache.sv:164:5
											wire [0:0] per_bank_core_rsp_idx;
											// Trace: src/VX_cache.sv:165:5
											wire [0:0] per_bank_core_rsp_ready;
											// Trace: src/VX_cache.sv:166:5
											wire [0:0] per_bank_mem_req_valid;
											// Trace: src/VX_cache.sv:167:5
											wire [25:0] per_bank_mem_req_addr;
											// Trace: src/VX_cache.sv:168:5
											wire [0:0] per_bank_mem_req_rw;
											// Trace: src/VX_cache.sv:169:5
											wire [63:0] per_bank_mem_req_byteen;
											// Trace: src/VX_cache.sv:170:5
											wire [511:0] per_bank_mem_req_data;
											// Trace: src/VX_cache.sv:171:5
											wire [4:0] per_bank_mem_req_tag;
											// Trace: src/VX_cache.sv:172:5
											wire [2:0] per_bank_mem_req_flags;
											// Trace: src/VX_cache.sv:173:5
											wire [0:0] per_bank_mem_req_ready;
											// Trace: src/VX_cache.sv:174:5
											wire [0:0] core_req_valid;
											// Trace: src/VX_cache.sv:175:5
											wire [27:0] core_req_addr;
											// Trace: src/VX_cache.sv:176:5
											wire [0:0] core_req_rw;
											// Trace: src/VX_cache.sv:177:5
											wire [15:0] core_req_byteen;
											// Trace: src/VX_cache.sv:178:5
											wire [127:0] core_req_data;
											// Trace: src/VX_cache.sv:179:5
											wire [2:0] core_req_tag;
											// Trace: src/VX_cache.sv:180:5
											wire [2:0] core_req_flags;
											// Trace: src/VX_cache.sv:181:5
											wire [0:0] core_req_ready;
											// Trace: src/VX_cache.sv:182:5
											wire [25:0] core_req_line_addr;
											// Trace: src/VX_cache.sv:183:5
											wire [0:0] core_req_bid;
											// Trace: src/VX_cache.sv:184:5
											wire [1:0] core_req_wsel;
											// Trace: src/VX_cache.sv:185:5
											wire [178:0] core_req_data_in;
											// Trace: src/VX_cache.sv:186:5
											wire [178:0] core_req_data_out;
											// Trace: src/VX_cache.sv:187:5
											genvar _gv_i_232;
											for (_gv_i_232 = 0; _gv_i_232 < NUM_REQS; _gv_i_232 = _gv_i_232 + 1) begin : g_core_req
												localparam i = _gv_i_232;
												// Trace: src/VX_cache.sv:188:9
												assign core_req_valid[i] = core_bus2_if[i].req_valid;
												// Trace: src/VX_cache.sv:189:9
												assign core_req_rw[i] = core_bus2_if[i].req_data[178];
												// Trace: src/VX_cache.sv:190:9
												assign core_req_byteen[i * 16+:16] = core_bus2_if[i].req_data[21-:16];
												// Trace: src/VX_cache.sv:191:9
												assign core_req_addr[i * 28+:28] = core_bus2_if[i].req_data[177-:28];
												// Trace: src/VX_cache.sv:192:9
												assign core_req_data[i * 128+:128] = core_bus2_if[i].req_data[149-:128];
												// Trace: src/VX_cache.sv:193:9
												assign core_req_tag[i * 3+:3] = core_bus2_if[i].req_data[2-:3];
												// Trace: src/VX_cache.sv:194:9
												assign core_req_flags[i * 3+:3] = sv2v_cast_3(core_bus2_if[i].req_data[5-:3]);
												// Trace: src/VX_cache.sv:195:9
												assign core_bus2_if[i].req_ready = core_req_ready[i];
											end
											// Trace: src/VX_cache.sv:197:5
											genvar _gv_i_233;
											for (_gv_i_233 = 0; _gv_i_233 < NUM_REQS; _gv_i_233 = _gv_i_233 + 1) begin : g_core_req_wsel
												localparam i = _gv_i_233;
												if (1) begin : g_wsel
													// Trace: src/VX_cache.sv:199:13
													assign core_req_wsel[i * 2+:2] = core_req_addr[i * 28+:WORD_SEL_BITS];
												end
											end
											// Trace: src/VX_cache.sv:204:5
											genvar _gv_i_234;
											for (_gv_i_234 = 0; _gv_i_234 < NUM_REQS; _gv_i_234 = _gv_i_234 + 1) begin : g_core_req_line_addr
												localparam i = _gv_i_234;
												// Trace: src/VX_cache.sv:205:9
												assign core_req_line_addr[i * 26+:26] = core_req_addr[(i * 28) + 2+:LINE_ADDR_WIDTH];
											end
											// Trace: src/VX_cache.sv:207:5
											genvar _gv_i_235;
											for (_gv_i_235 = 0; _gv_i_235 < NUM_REQS; _gv_i_235 = _gv_i_235 + 1) begin : g_core_req_bid
												localparam i = _gv_i_235;
												if (1) begin : g_singlebank
													// Trace: src/VX_cache.sv:211:13
													assign core_req_bid[i+:1] = 1'sb0;
												end
											end
											// Trace: src/VX_cache.sv:214:5
											genvar _gv_i_236;
											for (_gv_i_236 = 0; _gv_i_236 < NUM_REQS; _gv_i_236 = _gv_i_236 + 1) begin : g_core_req_data_in
												localparam i = _gv_i_236;
												// Trace: src/VX_cache.sv:215:9
												assign core_req_data_in[i * 179+:179] = {core_req_line_addr[i * 26+:26], core_req_rw[i], core_req_wsel[i * 2+:2], core_req_byteen[i * 16+:16], core_req_data[i * 128+:128], core_req_tag[i * 3+:3], core_req_flags[i * 3+:3]};
											end
											// Trace: src/VX_cache.sv:225:5
											assign per_bank_core_req_fire = per_bank_core_req_valid & per_bank_mem_req_ready;
											// Trace: src/VX_cache.sv:226:5
											localparam VX_gpu_pkg_PERF_CTR_BITS = 44;
											VX_stream_xbar #(
												.NUM_INPUTS(NUM_REQS),
												.NUM_OUTPUTS(NUM_BANKS),
												.DATAW(CORE_REQ_DATAW),
												.PERF_CTR_BITS(VX_gpu_pkg_PERF_CTR_BITS),
												.ARBITER("R"),
												.OUT_BUF(REQ_XBAR_BUF)
											) core_req_xbar(
												.clk(clk),
												.reset(reset),
												.collisions(),
												.valid_in(core_req_valid),
												.data_in(core_req_data_in),
												.sel_in(core_req_bid),
												.ready_in(core_req_ready),
												.valid_out(per_bank_core_req_valid),
												.data_out(core_req_data_out),
												.sel_out(per_bank_core_req_idx),
												.ready_out(per_bank_core_req_ready)
											);
											// Trace: src/VX_cache.sv:246:5
											genvar _gv_i_237;
											for (_gv_i_237 = 0; _gv_i_237 < NUM_BANKS; _gv_i_237 = _gv_i_237 + 1) begin : g_core_req_data_out
												localparam i = _gv_i_237;
												// Trace: src/VX_cache.sv:247:9
												assign {per_bank_core_req_addr[i * 26+:26], per_bank_core_req_rw[i], per_bank_core_req_wsel[i * 2+:2], per_bank_core_req_byteen[i * 16+:16], per_bank_core_req_data[i * 128+:128], per_bank_core_req_tag[i * 3+:3], per_bank_core_req_flags[i * 3+:3]} = core_req_data_out[i * 179+:179];
											end
											// Trace: src/VX_cache.sv:257:5
											genvar _gv_bank_id_1;
											for (_gv_bank_id_1 = 0; _gv_bank_id_1 < NUM_BANKS; _gv_bank_id_1 = _gv_bank_id_1 + 1) begin : g_banks
												localparam bank_id = _gv_bank_id_1;
												// Trace: src/VX_cache.sv:258:9
												VX_cache_bank #(
													.BANK_ID(bank_id),
													.INSTANCE_ID(""),
													.CACHE_SIZE(CACHE_SIZE),
													.LINE_SIZE(LINE_SIZE),
													.NUM_BANKS(NUM_BANKS),
													.NUM_WAYS(NUM_WAYS),
													.WORD_SIZE(WORD_SIZE),
													.NUM_REQS(NUM_REQS),
													.WRITE_ENABLE(WRITE_ENABLE),
													.WRITEBACK(WRITEBACK),
													.DIRTY_BYTES(DIRTY_BYTES),
													.REPL_POLICY(REPL_POLICY),
													.CRSQ_SIZE(CRSQ_SIZE),
													.MSHR_SIZE(MSHR_SIZE),
													.MREQ_SIZE(MREQ_SIZE),
													.TAG_WIDTH(TAG_WIDTH),
													.CORE_OUT_REG((CORE_RSP_BUF_ENABLE ? 0 : ((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : (CORE_OUT_BUF & 7) - 2))),
													.MEM_OUT_REG((MEM_REQ_BUF_ENABLE ? 0 : ((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : (MEM_OUT_BUF & 7) - 2)))
												) bank(
													.clk(clk),
													.reset(reset),
													.core_req_valid(per_bank_core_req_valid[bank_id]),
													.core_req_addr(per_bank_core_req_addr[bank_id * 26+:26]),
													.core_req_rw(per_bank_core_req_rw[bank_id]),
													.core_req_wsel(per_bank_core_req_wsel[bank_id * 2+:2]),
													.core_req_byteen(per_bank_core_req_byteen[bank_id * 16+:16]),
													.core_req_data(per_bank_core_req_data[bank_id * 128+:128]),
													.core_req_tag(per_bank_core_req_tag[bank_id * 3+:3]),
													.core_req_idx(per_bank_core_req_idx[bank_id+:1]),
													.core_req_flags(per_bank_core_req_flags[bank_id * 3+:3]),
													.core_req_ready(per_bank_core_req_ready[bank_id]),
													.core_rsp_valid(per_bank_core_rsp_valid[bank_id]),
													.core_rsp_data(per_bank_core_rsp_data[bank_id * 128+:128]),
													.core_rsp_tag(per_bank_core_rsp_tag[bank_id * 3+:3]),
													.core_rsp_idx(per_bank_core_rsp_idx[bank_id+:1]),
													.core_rsp_ready(per_bank_core_rsp_ready[bank_id]),
													.mem_req_valid(per_bank_mem_req_valid[bank_id]),
													.mem_req_addr(per_bank_mem_req_addr[bank_id * 26+:26]),
													.mem_req_rw(per_bank_mem_req_rw[bank_id]),
													.mem_req_byteen(per_bank_mem_req_byteen[bank_id * 64+:64]),
													.mem_req_data(per_bank_mem_req_data[bank_id * 512+:512]),
													.mem_req_tag(per_bank_mem_req_tag[bank_id * 5+:5]),
													.mem_req_flags(per_bank_mem_req_flags[bank_id * 3+:3]),
													.mem_req_ready(per_bank_mem_req_ready[bank_id]),
													.mem_rsp_valid(per_bank_mem_rsp_valid[bank_id]),
													.mem_rsp_data(per_bank_mem_rsp_data[bank_id * 512+:512]),
													.mem_rsp_tag(per_bank_mem_rsp_tag[bank_id * 5+:5]),
													.mem_rsp_ready(per_bank_mem_rsp_ready[bank_id]),
													.flush_begin(per_bank_flush_begin[bank_id]),
													.flush_uuid(flush_uuid),
													.flush_end(per_bank_flush_end[bank_id])
												);
											end
											// Trace: src/VX_cache.sv:312:5
											wire [130:0] core_rsp_data_in;
											// Trace: src/VX_cache.sv:313:5
											wire [130:0] core_rsp_data_out;
											// Trace: src/VX_cache.sv:314:5
											wire [0:0] core_rsp_valid_s;
											// Trace: src/VX_cache.sv:315:5
											wire [127:0] core_rsp_data_s;
											// Trace: src/VX_cache.sv:316:5
											wire [2:0] core_rsp_tag_s;
											// Trace: src/VX_cache.sv:317:5
											wire [0:0] core_rsp_ready_s;
											// Trace: src/VX_cache.sv:318:5
											genvar _gv_i_238;
											for (_gv_i_238 = 0; _gv_i_238 < NUM_BANKS; _gv_i_238 = _gv_i_238 + 1) begin : g_core_rsp_data_in
												localparam i = _gv_i_238;
												// Trace: src/VX_cache.sv:319:9
												assign core_rsp_data_in[i * 131+:131] = {per_bank_core_rsp_data[i * 128+:128], per_bank_core_rsp_tag[i * 3+:3]};
											end
											// Trace: src/VX_cache.sv:321:5
											VX_stream_xbar #(
												.NUM_INPUTS(NUM_BANKS),
												.NUM_OUTPUTS(NUM_REQS),
												.DATAW(CORE_RSP_DATAW),
												.ARBITER("R")
											) core_rsp_xbar(
												.clk(clk),
												.reset(reset),
												.collisions(),
												.valid_in(per_bank_core_rsp_valid),
												.data_in(core_rsp_data_in),
												.sel_in(per_bank_core_rsp_idx),
												.ready_in(per_bank_core_rsp_ready),
												.valid_out(core_rsp_valid_s),
												.data_out(core_rsp_data_out),
												.ready_out(core_rsp_ready_s),
												.sel_out()
											);
											// Trace: src/VX_cache.sv:339:5
											genvar _gv_i_239;
											for (_gv_i_239 = 0; _gv_i_239 < NUM_REQS; _gv_i_239 = _gv_i_239 + 1) begin : g_core_rsp_data_s
												localparam i = _gv_i_239;
												// Trace: src/VX_cache.sv:340:9
												assign {core_rsp_data_s[i * 128+:128], core_rsp_tag_s[i * 3+:3]} = core_rsp_data_out[i * 131+:131];
											end
											// Trace: src/VX_cache.sv:342:5
											genvar _gv_i_240;
											for (_gv_i_240 = 0; _gv_i_240 < NUM_REQS; _gv_i_240 = _gv_i_240 + 1) begin : g_core_rsp_buf
												localparam i = _gv_i_240;
												// Trace: src/VX_cache.sv:343:9
												VX_elastic_buffer #(
													.DATAW(131),
													.SIZE((CORE_RSP_BUF_ENABLE ? ((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : 2) : 0)),
													.OUT_REG(((CORE_OUT_BUF & 7) < 2 ? CORE_OUT_BUF & 7 : (CORE_OUT_BUF & 7) - 2))
												) core_rsp_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(core_rsp_valid_s[i]),
													.ready_in(core_rsp_ready_s[i]),
													.data_in({core_rsp_data_s[i * 128+:128], core_rsp_tag_s[i * 3+:3]}),
													.data_out({core_bus2_if[i].rsp_data[130-:128], core_bus2_if[i].rsp_data[2-:3]}),
													.valid_out(core_bus2_if[i].rsp_valid),
													.ready_out(core_bus2_if[i].rsp_ready)
												);
											end
											// Trace: src/VX_cache.sv:358:5
											wire [610:0] per_bank_mem_req_pdata;
											// Trace: src/VX_cache.sv:359:5
											genvar _gv_i_241;
											for (_gv_i_241 = 0; _gv_i_241 < NUM_BANKS; _gv_i_241 = _gv_i_241 + 1) begin : g_per_bank_mem_req_pdata
												localparam i = _gv_i_241;
												// Trace: src/VX_cache.sv:360:9
												assign per_bank_mem_req_pdata[i * 611+:611] = {per_bank_mem_req_rw[i], per_bank_mem_req_addr[i * 26+:26], per_bank_mem_req_data[i * 512+:512], per_bank_mem_req_byteen[i * 64+:64], per_bank_mem_req_flags[i * 3+:3], per_bank_mem_req_tag[i * 5+:5]};
											end
											// Trace: src/VX_cache.sv:369:5
											wire [0:0] mem_req_valid;
											// Trace: src/VX_cache.sv:370:5
											wire [610:0] mem_req_pdata;
											// Trace: src/VX_cache.sv:371:5
											wire [0:0] mem_req_ready;
											// Trace: src/VX_cache.sv:372:5
											wire [0:0] mem_req_sel_out;
											// Trace: src/VX_cache.sv:373:5
											VX_stream_arb #(
												.NUM_INPUTS(NUM_BANKS),
												.NUM_OUTPUTS(MEM_PORTS),
												.DATAW(MEM_REQ_DATAW),
												.ARBITER("R")
											) mem_req_arb(
												.clk(clk),
												.reset(reset),
												.valid_in(per_bank_mem_req_valid),
												.data_in(per_bank_mem_req_pdata),
												.ready_in(per_bank_mem_req_ready),
												.valid_out(mem_req_valid),
												.data_out(mem_req_pdata),
												.ready_out(mem_req_ready),
												.sel_out(mem_req_sel_out)
											);
											// Trace: src/VX_cache.sv:389:5
											genvar _gv_i_242;
											for (_gv_i_242 = 0; _gv_i_242 < MEM_PORTS; _gv_i_242 = _gv_i_242 + 1) begin : g_mem_req_buf
												localparam i = _gv_i_242;
												// Trace: src/VX_cache.sv:390:9
												wire mem_req_rw;
												// Trace: src/VX_cache.sv:391:9
												wire [25:0] mem_req_addr;
												// Trace: src/VX_cache.sv:392:9
												wire [511:0] mem_req_data;
												// Trace: src/VX_cache.sv:393:9
												wire [63:0] mem_req_byteen;
												// Trace: src/VX_cache.sv:394:9
												wire [2:0] mem_req_flags;
												// Trace: src/VX_cache.sv:395:9
												wire [4:0] mem_req_tag;
												// Trace: src/VX_cache.sv:396:9
												assign {mem_req_rw, mem_req_addr, mem_req_data, mem_req_byteen, mem_req_flags, mem_req_tag} = mem_req_pdata[i * 611+:611];
												// Trace: src/VX_cache.sv:404:9
												wire [25:0] mem_req_addr_w;
												// Trace: src/VX_cache.sv:405:9
												wire [4:0] mem_req_tag_w;
												// Trace: src/VX_cache.sv:406:9
												wire [2:0] mem_req_flags_w;
												if (1) begin : g_mem_req_tag
													// Trace: src/VX_cache.sv:425:13
													assign mem_req_addr_w = mem_req_addr;
													// Trace: src/VX_cache.sv:426:13
													assign mem_req_tag_w = mem_req_tag;
												end
												// Trace: src/VX_cache.sv:428:9
												VX_elastic_buffer #(
													.DATAW(611),
													.SIZE((MEM_REQ_BUF_ENABLE ? ((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : 2) : 0)),
													.OUT_REG(((MEM_OUT_BUF & 7) < 2 ? MEM_OUT_BUF & 7 : (MEM_OUT_BUF & 7) - 2))
												) mem_req_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(mem_req_valid[i]),
													.ready_in(mem_req_ready[i]),
													.data_in({mem_req_rw, mem_req_byteen, mem_req_addr_w, mem_req_data, mem_req_tag_w, mem_req_flags}),
													.data_out({mem_bus_tmp_if[i].req_data[610], mem_bus_tmp_if[i].req_data[71-:64], mem_bus_tmp_if[i].req_data[609-:26], mem_bus_tmp_if[i].req_data[583-:512], mem_bus_tmp_if[i].req_data[4-:5], mem_req_flags_w}),
													.valid_out(mem_bus_tmp_if[i].req_valid),
													.ready_out(mem_bus_tmp_if[i].req_ready)
												);
												if (1) begin : g_mem_req_flags
													// Trace: src/VX_cache.sv:443:13
													assign mem_bus_tmp_if[i].req_data[7-:3] = mem_req_flags_w;
												end
												if (WRITE_ENABLE) begin : g_mem_bus_if
													// Trace: src/VX_cache.sv:448:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
													// Trace: src/VX_cache.sv:449:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[i].req_data;
													// Trace: src/VX_cache.sv:450:5
													assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_ready;
													// Trace: src/VX_cache.sv:451:5
													assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_valid;
													// Trace: src/VX_cache.sv:452:5
													assign mem_bus_tmp_if[i].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_data;
													// Trace: src/VX_cache.sv:453:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
												end
												else begin : g_mem_bus_if_ro
													// Trace: src/VX_cache.sv:455:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[i].req_valid;
													// Trace: src/VX_cache.sv:456:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[610] = 0;
													// Trace: src/VX_cache.sv:457:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[609-:26] = mem_bus_tmp_if[i].req_data[609-:26];
													// Trace: src/VX_cache.sv:458:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[583-:512] = 1'sb0;
													// Trace: src/VX_cache.sv:459:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[71-:64] = 1'sb1;
													// Trace: src/VX_cache.sv:460:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[7-:3] = mem_bus_tmp_if[i].req_data[7-:3];
													// Trace: src/VX_cache.sv:461:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_data[4-:5] = mem_bus_tmp_if[i].req_data[4-:5];
													// Trace: src/VX_cache.sv:462:5
													assign mem_bus_tmp_if[i].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].req_ready;
													// Trace: src/VX_cache.sv:463:5
													assign mem_bus_tmp_if[i].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_valid;
													// Trace: src/VX_cache.sv:464:5
													assign mem_bus_tmp_if[i].rsp_data[516-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_data[516-:512];
													// Trace: src/VX_cache.sv:465:5
													assign mem_bus_tmp_if[i].rsp_data[4-:5] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_data[4-:5];
													// Trace: src/VX_cache.sv:466:5
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_cache_wrap[_gv_i_192].cache_wrap.mem_bus_cache_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[i].rsp_ready;
												end
											end
										end
										assign cache.clk = clk;
										assign cache.reset = reset;
									end
								end
								assign cache_wrap.clk = clk;
								assign cache_wrap.reset = reset;
							end
							// Trace: src/VX_cache_cluster.sv:120:5
							genvar _gv_i_193;
							for (_gv_i_193 = 0; _gv_i_193 < MEM_PORTS; _gv_i_193 = _gv_i_193 + 1) begin : g_mem_bus_if
								localparam i = _gv_i_193;
								// Trace: src/VX_cache_cluster.sv:121:9
								// expanded interface instance: arb_core_bus_tmp_if
								localparam _param_E788B_DATA_SIZE = LINE_SIZE;
								localparam _param_E788B_TAG_WIDTH = MEM_TAG_WIDTH;
								genvar _arr_E788B;
								for (_arr_E788B = 0; _arr_E788B <= 0; _arr_E788B = _arr_E788B + 1) begin : arb_core_bus_tmp_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_E788B_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_E788B_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:8:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:12:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:20:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:24:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire [611:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire [517:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:30:5
									// Trace: src/VX_mem_bus_if.sv:38:5
								end
								// Trace: src/VX_cache_cluster.sv:125:9
								// expanded interface instance: mem_bus_tmp_if
								localparam _param_4FE36_DATA_SIZE = LINE_SIZE;
								localparam _param_4FE36_TAG_WIDTH = MEM_TAG_WIDTH + 0;
								genvar _arr_4FE36;
								for (_arr_4FE36 = 0; _arr_4FE36 <= 0; _arr_4FE36 = _arr_4FE36 + 1) begin : mem_bus_tmp_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_4FE36_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_4FE36_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:8:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:12:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:20:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:24:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire [611:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire [517:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:30:5
									// Trace: src/VX_mem_bus_if.sv:38:5
								end
								genvar _gv_j_20;
								for (_gv_j_20 = 0; _gv_j_20 < NUM_CACHES; _gv_j_20 = _gv_j_20 + 1) begin : g_arb_core_bus_tmp_if
									localparam j = _gv_j_20;
									// Trace: src/VX_cache_cluster.sv:130:5
									assign arb_core_bus_tmp_if[j].req_valid = cache_mem_bus_if[(j * MEM_PORTS) + i].req_valid;
									// Trace: src/VX_cache_cluster.sv:131:5
									assign arb_core_bus_tmp_if[j].req_data = cache_mem_bus_if[(j * MEM_PORTS) + i].req_data;
									// Trace: src/VX_cache_cluster.sv:132:5
									assign cache_mem_bus_if[(j * MEM_PORTS) + i].req_ready = arb_core_bus_tmp_if[j].req_ready;
									// Trace: src/VX_cache_cluster.sv:133:5
									assign cache_mem_bus_if[(j * MEM_PORTS) + i].rsp_valid = arb_core_bus_tmp_if[j].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:134:5
									assign cache_mem_bus_if[(j * MEM_PORTS) + i].rsp_data = arb_core_bus_tmp_if[j].rsp_data;
									// Trace: src/VX_cache_cluster.sv:135:5
									assign arb_core_bus_tmp_if[j].rsp_ready = cache_mem_bus_if[(j * MEM_PORTS) + i].rsp_ready;
								end
								// Trace: src/VX_cache_cluster.sv:137:9
								// expanded module instance: mem_arb
								localparam _bbase_7277A_bus_in_if = 0;
								localparam _bbase_7277A_bus_out_if = 0;
								localparam _param_7277A_NUM_INPUTS = NUM_CACHES;
								localparam _param_7277A_NUM_OUTPUTS = 1;
								localparam _param_7277A_DATA_SIZE = LINE_SIZE;
								localparam _param_7277A_TAG_WIDTH = MEM_TAG_WIDTH;
								localparam _param_7277A_TAG_SEL_IDX = TAG_SEL_IDX;
								localparam _param_7277A_ARBITER = "R";
								localparam _param_7277A_REQ_OUT_BUF = 0;
								localparam _param_7277A_RSP_OUT_BUF = 0;
								if (1) begin : mem_arb
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_arb.sv:2:15
									localparam NUM_INPUTS = _param_7277A_NUM_INPUTS;
									// Trace: src/VX_mem_arb.sv:3:15
									localparam NUM_OUTPUTS = _param_7277A_NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:4:15
									localparam DATA_SIZE = _param_7277A_DATA_SIZE;
									// Trace: src/VX_mem_arb.sv:5:15
									localparam TAG_WIDTH = _param_7277A_TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:6:15
									localparam TAG_SEL_IDX = _param_7277A_TAG_SEL_IDX;
									// Trace: src/VX_mem_arb.sv:7:15
									localparam REQ_OUT_BUF = _param_7277A_REQ_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:8:15
									localparam RSP_OUT_BUF = _param_7277A_RSP_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:9:15
									localparam ARBITER = _param_7277A_ARBITER;
									// Trace: src/VX_mem_arb.sv:10:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_arb.sv:11:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_arb.sv:12:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_arb.sv:14:5
									wire clk;
									// Trace: src/VX_mem_arb.sv:15:5
									wire reset;
									// Trace: src/VX_mem_arb.sv:16:5
									localparam _mbase_bus_in_if = 0;
									// Trace: src/VX_mem_arb.sv:17:5
									localparam _mbase_bus_out_if = 0;
									// Trace: src/VX_mem_arb.sv:19:5
									localparam DATA_WIDTH = 512;
									// Trace: src/VX_mem_arb.sv:20:5
									localparam LOG_NUM_REQS = 0;
									// Trace: src/VX_mem_arb.sv:21:5
									localparam REQ_DATAW = 606 + TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:22:5
									localparam RSP_DATAW = DATA_WIDTH + TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:23:5
									localparam SEL_COUNT = NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:24:5
									wire [0:0] req_valid_in;
									// Trace: src/VX_mem_arb.sv:25:5
									wire [REQ_DATAW - 1:0] req_data_in;
									// Trace: src/VX_mem_arb.sv:26:5
									wire [0:0] req_ready_in;
									// Trace: src/VX_mem_arb.sv:27:5
									wire [0:0] req_valid_out;
									// Trace: src/VX_mem_arb.sv:28:5
									wire [REQ_DATAW - 1:0] req_data_out;
									// Trace: src/VX_mem_arb.sv:29:5
									wire [0:0] req_sel_out;
									// Trace: src/VX_mem_arb.sv:30:5
									wire [0:0] req_ready_out;
									// Trace: src/VX_mem_arb.sv:31:5
									genvar _gv_i_183;
									for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
										localparam i = _gv_i_183;
										// Trace: src/VX_mem_arb.sv:32:9
										assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].arb_core_bus_tmp_if[i + _mbase_bus_in_if].req_valid;
										// Trace: src/VX_mem_arb.sv:33:9
										assign req_data_in[i * 612+:612] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].arb_core_bus_tmp_if[i + _mbase_bus_in_if].req_data;
										// Trace: src/VX_mem_arb.sv:34:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].arb_core_bus_tmp_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:36:5
									VX_stream_arb #(
										.NUM_INPUTS(NUM_INPUTS),
										.NUM_OUTPUTS(NUM_OUTPUTS),
										.DATAW(REQ_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(REQ_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(req_valid_in),
										.ready_in(req_ready_in),
										.data_in(req_data_in),
										.data_out(req_data_out),
										.sel_out(req_sel_out),
										.valid_out(req_valid_out),
										.ready_out(req_ready_out)
									);
									// Trace: src/VX_mem_arb.sv:53:5
									genvar _gv_i_184;
									for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
										localparam i = _gv_i_184;
										// Trace: src/VX_mem_arb.sv:54:9
										wire [TAG_WIDTH - 1:0] req_tag_out;
										// Trace: src/VX_mem_arb.sv:55:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
										// Trace: src/VX_mem_arb.sv:56:9
										assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[611], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[610-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[584-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[72-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[8-:3], req_tag_out} = req_data_out[i * 612+:612];
										// Trace: src/VX_mem_arb.sv:64:9
										assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_ready;
										if (1) begin : g_req_tag_out
											// Trace: src/VX_mem_arb.sv:76:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].req_data[5-:6] = req_tag_out;
										end
									end
									// Trace: src/VX_mem_arb.sv:79:5
									wire [0:0] rsp_valid_out;
									// Trace: src/VX_mem_arb.sv:80:5
									wire [RSP_DATAW - 1:0] rsp_data_out;
									// Trace: src/VX_mem_arb.sv:81:5
									wire [0:0] rsp_ready_out;
									// Trace: src/VX_mem_arb.sv:82:5
									wire [0:0] rsp_valid_in;
									// Trace: src/VX_mem_arb.sv:83:5
									wire [RSP_DATAW - 1:0] rsp_data_in;
									// Trace: src/VX_mem_arb.sv:84:5
									wire [0:0] rsp_ready_in;
									// Trace: src/VX_mem_arb.sv:85:5
									if (1) begin : g_rsp_arb
										genvar _gv_i_186;
										for (_gv_i_186 = 0; _gv_i_186 < NUM_OUTPUTS; _gv_i_186 = _gv_i_186 + 1) begin : g_rsp_data_in
											localparam i = _gv_i_186;
											// Trace: src/VX_mem_arb.sv:120:13
											assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_valid;
											// Trace: src/VX_mem_arb.sv:121:13
											assign rsp_data_in[i * 518+:518] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_data;
											// Trace: src/VX_mem_arb.sv:122:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].mem_bus_tmp_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
										end
										// Trace: src/VX_mem_arb.sv:124:9
										VX_stream_arb #(
											.NUM_INPUTS(NUM_OUTPUTS),
											.NUM_OUTPUTS(NUM_INPUTS),
											.DATAW(RSP_DATAW),
											.ARBITER(ARBITER),
											.OUT_BUF(RSP_OUT_BUF)
										) req_arb(
											.clk(clk),
											.reset(reset),
											.valid_in(rsp_valid_in),
											.ready_in(rsp_ready_in),
											.data_in(rsp_data_in),
											.data_out(rsp_data_out),
											.valid_out(rsp_valid_out),
											.ready_out(rsp_ready_out),
											.sel_out()
										);
									end
									// Trace: src/VX_mem_arb.sv:142:5
									genvar _gv_i_187;
									for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
										localparam i = _gv_i_187;
										// Trace: src/VX_mem_arb.sv:143:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].arb_core_bus_tmp_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
										// Trace: src/VX_mem_arb.sv:144:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].arb_core_bus_tmp_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 518+:518];
										// Trace: src/VX_mem_arb.sv:145:9
										assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache.g_mem_bus_if[_gv_i_193].arb_core_bus_tmp_if[i + _mbase_bus_in_if].rsp_ready;
									end
								end
								assign mem_arb.clk = clk;
								assign mem_arb.reset = reset;
								if (WRITE_ENABLE) begin : g_we
									// Trace: src/VX_cache_cluster.sv:153:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[0].req_valid;
									// Trace: src/VX_cache_cluster.sv:154:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data = mem_bus_tmp_if[0].req_data;
									// Trace: src/VX_cache_cluster.sv:155:5
									assign mem_bus_tmp_if[0].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
									// Trace: src/VX_cache_cluster.sv:156:5
									assign mem_bus_tmp_if[0].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:157:5
									assign mem_bus_tmp_if[0].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
									// Trace: src/VX_cache_cluster.sv:158:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[0].rsp_ready;
								end
								else begin : g_ro
									// Trace: src/VX_cache_cluster.sv:160:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_valid = mem_bus_tmp_if[0].req_valid;
									// Trace: src/VX_cache_cluster.sv:161:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data[611] = 0;
									// Trace: src/VX_cache_cluster.sv:162:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data[610-:26] = mem_bus_tmp_if[0].req_data[610-:26];
									// Trace: src/VX_cache_cluster.sv:163:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data[584-:512] = 1'sb0;
									// Trace: src/VX_cache_cluster.sv:164:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data[72-:64] = 1'sb1;
									// Trace: src/VX_cache_cluster.sv:165:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data[8-:3] = mem_bus_tmp_if[0].req_data[8-:3];
									// Trace: src/VX_cache_cluster.sv:166:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_data[5-:6] = mem_bus_tmp_if[0].req_data[5-:6];
									// Trace: src/VX_cache_cluster.sv:167:5
									assign mem_bus_tmp_if[0].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
									// Trace: src/VX_cache_cluster.sv:168:5
									assign mem_bus_tmp_if[0].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
									// Trace: src/VX_cache_cluster.sv:169:5
									assign mem_bus_tmp_if[0].rsp_data[517-:512] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[517-:512];
									// Trace: src/VX_cache_cluster.sv:170:5
									assign mem_bus_tmp_if[0].rsp_data[5-:6] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_data[5-:6];
									// Trace: src/VX_cache_cluster.sv:171:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.dcache_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = mem_bus_tmp_if[0].rsp_ready;
								end
							end
						end
						assign dcache.clk = clk;
						assign dcache.reset = dcache_reset;
						// Trace: src/VX_socket.sv:97:5
						genvar _gv_i_180;
						localparam VX_gpu_pkg_L1_MEM_TAG_WIDTH = VX_gpu_pkg_DCACHE_MEM_TAG_WIDTH;
						localparam VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH = 7;
						for (_gv_i_180 = 0; _gv_i_180 < VX_gpu_pkg_DCACHE_NUM_REQS; _gv_i_180 = _gv_i_180 + 1) begin : g_mem_bus_if
							localparam i = _gv_i_180;
							if (i == 0) begin : g_i0
								// Trace: src/VX_socket.sv:99:13
								// expanded interface instance: l1_mem_bus_if
								localparam _param_70CB9_DATA_SIZE = 64;
								localparam _param_70CB9_TAG_WIDTH = VX_gpu_pkg_L1_MEM_TAG_WIDTH;
								genvar _arr_70CB9;
								for (_arr_70CB9 = 0; _arr_70CB9 <= 1; _arr_70CB9 = _arr_70CB9 + 1) begin : l1_mem_bus_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_70CB9_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_70CB9_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:8:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:12:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:20:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:24:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire [611:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire [517:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:30:5
									// Trace: src/VX_mem_bus_if.sv:38:5
								end
								// Trace: src/VX_socket.sv:103:13
								// expanded interface instance: l1_mem_arb_bus_if
								localparam _param_D5D25_DATA_SIZE = 64;
								localparam _param_D5D25_TAG_WIDTH = VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH;
								genvar _arr_D5D25;
								for (_arr_D5D25 = 0; _arr_D5D25 <= 0; _arr_D5D25 = _arr_D5D25 + 1) begin : l1_mem_arb_bus_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_D5D25_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_D5D25_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:8:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:12:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:20:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:24:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire [612:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire [518:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:30:5
									// Trace: src/VX_mem_bus_if.sv:38:5
								end
								// Trace: src/VX_socket.sv:108:5
								assign l1_mem_bus_if[0].req_valid = icache_mem_bus_if[0].req_valid;
								// Trace: src/VX_socket.sv:109:5
								assign l1_mem_bus_if[0].req_data[611] = icache_mem_bus_if[0].req_data[610];
								// Trace: src/VX_socket.sv:110:5
								assign l1_mem_bus_if[0].req_data[610-:26] = icache_mem_bus_if[0].req_data[609-:26];
								// Trace: src/VX_socket.sv:111:5
								assign l1_mem_bus_if[0].req_data[584-:512] = icache_mem_bus_if[0].req_data[583-:512];
								// Trace: src/VX_socket.sv:112:5
								assign l1_mem_bus_if[0].req_data[72-:64] = icache_mem_bus_if[0].req_data[71-:64];
								// Trace: src/VX_socket.sv:113:5
								assign l1_mem_bus_if[0].req_data[8-:3] = icache_mem_bus_if[0].req_data[7-:3];
								if (1) begin : genblk1
									if (1) begin : genblk1
										if (1) begin : genblk1
											// Trace: src/VX_socket.sv:117:17
											assign l1_mem_bus_if[0].req_data[5-:6] = {icache_mem_bus_if[0].req_data[4-:1], 1'b0, icache_mem_bus_if[0].req_data[3-:4]};
										end
									end
								end
								// Trace: src/VX_socket.sv:131:5
								assign icache_mem_bus_if[0].req_ready = l1_mem_bus_if[0].req_ready;
								// Trace: src/VX_socket.sv:132:5
								assign icache_mem_bus_if[0].rsp_valid = l1_mem_bus_if[0].rsp_valid;
								// Trace: src/VX_socket.sv:133:5
								assign icache_mem_bus_if[0].rsp_data[516-:512] = l1_mem_bus_if[0].rsp_data[517-:512];
								if (1) begin : genblk2
									if (1) begin : genblk1
										if (1) begin : genblk1
											// Trace: src/VX_socket.sv:137:17
											assign icache_mem_bus_if[0].rsp_data[4-:5] = {l1_mem_bus_if[0].rsp_data[5-:1], l1_mem_bus_if[0].rsp_data[3:0]};
										end
									end
								end
								// Trace: src/VX_socket.sv:151:5
								assign l1_mem_bus_if[0].rsp_ready = icache_mem_bus_if[0].rsp_ready;
								// Trace: src/VX_socket.sv:154:5
								assign l1_mem_bus_if[1].req_valid = dcache_mem_bus_if[0].req_valid;
								// Trace: src/VX_socket.sv:155:5
								assign l1_mem_bus_if[1].req_data[611] = dcache_mem_bus_if[0].req_data[611];
								// Trace: src/VX_socket.sv:156:5
								assign l1_mem_bus_if[1].req_data[610-:26] = dcache_mem_bus_if[0].req_data[610-:26];
								// Trace: src/VX_socket.sv:157:5
								assign l1_mem_bus_if[1].req_data[584-:512] = dcache_mem_bus_if[0].req_data[584-:512];
								// Trace: src/VX_socket.sv:158:5
								assign l1_mem_bus_if[1].req_data[72-:64] = dcache_mem_bus_if[0].req_data[72-:64];
								// Trace: src/VX_socket.sv:159:5
								assign l1_mem_bus_if[1].req_data[8-:3] = dcache_mem_bus_if[0].req_data[8-:3];
								if (1) begin : genblk3
									// Trace: src/VX_socket.sv:175:9
									assign l1_mem_bus_if[1].req_data[5-:6] = dcache_mem_bus_if[0].req_data[5-:6];
								end
								// Trace: src/VX_socket.sv:177:5
								assign dcache_mem_bus_if[0].req_ready = l1_mem_bus_if[1].req_ready;
								// Trace: src/VX_socket.sv:178:5
								assign dcache_mem_bus_if[0].rsp_valid = l1_mem_bus_if[1].rsp_valid;
								// Trace: src/VX_socket.sv:179:5
								assign dcache_mem_bus_if[0].rsp_data[517-:512] = l1_mem_bus_if[1].rsp_data[517-:512];
								if (1) begin : genblk4
									// Trace: src/VX_socket.sv:195:9
									assign dcache_mem_bus_if[0].rsp_data[5-:6] = l1_mem_bus_if[1].rsp_data[5-:6];
								end
								// Trace: src/VX_socket.sv:197:5
								assign l1_mem_bus_if[1].rsp_ready = dcache_mem_bus_if[0].rsp_ready;
								// Trace: src/VX_socket.sv:199:13
								// expanded module instance: mem_arb
								localparam _bbase_7277A_bus_in_if = 0;
								localparam _bbase_7277A_bus_out_if = 0;
								localparam _param_7277A_NUM_INPUTS = 2;
								localparam _param_7277A_NUM_OUTPUTS = 1;
								localparam _param_7277A_DATA_SIZE = 64;
								localparam _param_7277A_TAG_WIDTH = VX_gpu_pkg_L1_MEM_TAG_WIDTH;
								localparam _param_7277A_TAG_SEL_IDX = 0;
								localparam _param_7277A_ARBITER = "P";
								localparam _param_7277A_REQ_OUT_BUF = 3;
								localparam _param_7277A_RSP_OUT_BUF = 3;
								if (1) begin : mem_arb
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_arb.sv:2:15
									localparam NUM_INPUTS = _param_7277A_NUM_INPUTS;
									// Trace: src/VX_mem_arb.sv:3:15
									localparam NUM_OUTPUTS = _param_7277A_NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:4:15
									localparam DATA_SIZE = _param_7277A_DATA_SIZE;
									// Trace: src/VX_mem_arb.sv:5:15
									localparam TAG_WIDTH = _param_7277A_TAG_WIDTH;
									// Trace: src/VX_mem_arb.sv:6:15
									localparam TAG_SEL_IDX = _param_7277A_TAG_SEL_IDX;
									// Trace: src/VX_mem_arb.sv:7:15
									localparam REQ_OUT_BUF = _param_7277A_REQ_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:8:15
									localparam RSP_OUT_BUF = _param_7277A_RSP_OUT_BUF;
									// Trace: src/VX_mem_arb.sv:9:15
									localparam ARBITER = _param_7277A_ARBITER;
									// Trace: src/VX_mem_arb.sv:10:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_arb.sv:11:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_arb.sv:12:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_arb.sv:14:5
									wire clk;
									// Trace: src/VX_mem_arb.sv:15:5
									wire reset;
									// Trace: src/VX_mem_arb.sv:16:5
									localparam _mbase_bus_in_if = 0;
									// Trace: src/VX_mem_arb.sv:17:5
									localparam _mbase_bus_out_if = 0;
									// Trace: src/VX_mem_arb.sv:19:5
									localparam DATA_WIDTH = 512;
									// Trace: src/VX_mem_arb.sv:20:5
									localparam LOG_NUM_REQS = 1;
									// Trace: src/VX_mem_arb.sv:21:5
									localparam REQ_DATAW = 612;
									// Trace: src/VX_mem_arb.sv:22:5
									localparam RSP_DATAW = 518;
									// Trace: src/VX_mem_arb.sv:23:5
									localparam SEL_COUNT = NUM_OUTPUTS;
									// Trace: src/VX_mem_arb.sv:24:5
									wire [1:0] req_valid_in;
									// Trace: src/VX_mem_arb.sv:25:5
									wire [1223:0] req_data_in;
									// Trace: src/VX_mem_arb.sv:26:5
									wire [1:0] req_ready_in;
									// Trace: src/VX_mem_arb.sv:27:5
									wire [0:0] req_valid_out;
									// Trace: src/VX_mem_arb.sv:28:5
									wire [611:0] req_data_out;
									// Trace: src/VX_mem_arb.sv:29:5
									wire [0:0] req_sel_out;
									// Trace: src/VX_mem_arb.sv:30:5
									wire [0:0] req_ready_out;
									// Trace: src/VX_mem_arb.sv:31:5
									genvar _gv_i_183;
									for (_gv_i_183 = 0; _gv_i_183 < NUM_INPUTS; _gv_i_183 = _gv_i_183 + 1) begin : g_req_data_in
										localparam i = _gv_i_183;
										// Trace: src/VX_mem_arb.sv:32:9
										assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_bus_if[i + _mbase_bus_in_if].req_valid;
										// Trace: src/VX_mem_arb.sv:33:9
										assign req_data_in[i * 612+:612] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_bus_if[i + _mbase_bus_in_if].req_data;
										// Trace: src/VX_mem_arb.sv:34:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_bus_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
									end
									// Trace: src/VX_mem_arb.sv:36:5
									VX_stream_arb #(
										.NUM_INPUTS(NUM_INPUTS),
										.NUM_OUTPUTS(NUM_OUTPUTS),
										.DATAW(REQ_DATAW),
										.ARBITER(ARBITER),
										.OUT_BUF(REQ_OUT_BUF)
									) req_arb(
										.clk(clk),
										.reset(reset),
										.valid_in(req_valid_in),
										.ready_in(req_ready_in),
										.data_in(req_data_in),
										.data_out(req_data_out),
										.sel_out(req_sel_out),
										.valid_out(req_valid_out),
										.ready_out(req_ready_out)
									);
									// Trace: src/VX_mem_arb.sv:53:5
									genvar _gv_i_184;
									for (_gv_i_184 = 0; _gv_i_184 < NUM_OUTPUTS; _gv_i_184 = _gv_i_184 + 1) begin : g_bus_out_if
										localparam i = _gv_i_184;
										// Trace: src/VX_mem_arb.sv:54:9
										wire [5:0] req_tag_out;
										// Trace: src/VX_mem_arb.sv:55:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
										// Trace: src/VX_mem_arb.sv:56:9
										assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_data[612], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_data[611-:26], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_data[585-:512], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_data[73-:64], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_data[9-:3], req_tag_out} = req_data_out[i * 612+:612];
										// Trace: src/VX_mem_arb.sv:64:9
										assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_ready;
										if (1) begin : g_req_tag_sel_out
											// Trace: src/VX_mem_arb.sv:66:13
											VX_bits_insert #(
												.N(TAG_WIDTH),
												.S(LOG_NUM_REQS),
												.POS(TAG_SEL_IDX)
											) bits_insert(
												.data_in(req_tag_out),
												.ins_in(req_sel_out[i+:1]),
												.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].req_data[6-:7])
											);
										end
									end
									// Trace: src/VX_mem_arb.sv:79:5
									wire [1:0] rsp_valid_out;
									// Trace: src/VX_mem_arb.sv:80:5
									wire [1035:0] rsp_data_out;
									// Trace: src/VX_mem_arb.sv:81:5
									wire [1:0] rsp_ready_out;
									// Trace: src/VX_mem_arb.sv:82:5
									wire [0:0] rsp_valid_in;
									// Trace: src/VX_mem_arb.sv:83:5
									wire [517:0] rsp_data_in;
									// Trace: src/VX_mem_arb.sv:84:5
									wire [0:0] rsp_ready_in;
									// Trace: src/VX_mem_arb.sv:85:5
									if (1) begin : g_rsp_select
										// Trace: src/VX_mem_arb.sv:86:9
										wire [0:0] rsp_sel_in;
										genvar _gv_i_185;
										for (_gv_i_185 = 0; _gv_i_185 < NUM_OUTPUTS; _gv_i_185 = _gv_i_185 + 1) begin : g_rsp_data_in
											localparam i = _gv_i_185;
											// Trace: src/VX_mem_arb.sv:88:13
											wire [5:0] rsp_tag_out;
											// Trace: src/VX_mem_arb.sv:89:13
											VX_bits_remove #(
												.N(7),
												.S(LOG_NUM_REQS),
												.POS(TAG_SEL_IDX)
											) bits_remove(
												.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].rsp_data[6-:7]),
												.sel_out(rsp_sel_in[i+:1]),
												.data_out(rsp_tag_out)
											);
											// Trace: src/VX_mem_arb.sv:98:13
											assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].rsp_valid;
											// Trace: src/VX_mem_arb.sv:99:13
											assign rsp_data_in[i * 518+:518] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].rsp_data[518-:512], rsp_tag_out};
											// Trace: src/VX_mem_arb.sv:100:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_arb_bus_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
										end
										// Trace: src/VX_mem_arb.sv:102:9
										VX_stream_switch #(
											.NUM_INPUTS(NUM_OUTPUTS),
											.NUM_OUTPUTS(NUM_INPUTS),
											.DATAW(RSP_DATAW),
											.OUT_BUF(RSP_OUT_BUF)
										) rsp_switch(
											.clk(clk),
											.reset(reset),
											.sel_in(rsp_sel_in),
											.valid_in(rsp_valid_in),
											.ready_in(rsp_ready_in),
											.data_in(rsp_data_in),
											.data_out(rsp_data_out),
											.valid_out(rsp_valid_out),
											.ready_out(rsp_ready_out)
										);
									end
									// Trace: src/VX_mem_arb.sv:142:5
									genvar _gv_i_187;
									for (_gv_i_187 = 0; _gv_i_187 < NUM_INPUTS; _gv_i_187 = _gv_i_187 + 1) begin : g_output
										localparam i = _gv_i_187;
										// Trace: src/VX_mem_arb.sv:143:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_bus_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
										// Trace: src/VX_mem_arb.sv:144:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_bus_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 518+:518];
										// Trace: src/VX_mem_arb.sv:145:9
										assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_mem_bus_if[_gv_i_180].g_i0.l1_mem_bus_if[i + _mbase_bus_in_if].rsp_ready;
									end
								end
								assign mem_arb.clk = clk;
								assign mem_arb.reset = reset;
								// Trace: src/VX_socket.sv:214:5
								assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[0 + _mbase_mem_bus_if].req_valid = l1_mem_arb_bus_if[0].req_valid;
								// Trace: src/VX_socket.sv:215:5
								assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[0 + _mbase_mem_bus_if].req_data = l1_mem_arb_bus_if[0].req_data;
								// Trace: src/VX_socket.sv:216:5
								assign l1_mem_arb_bus_if[0].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[0 + _mbase_mem_bus_if].req_ready;
								// Trace: src/VX_socket.sv:217:5
								assign l1_mem_arb_bus_if[0].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[0 + _mbase_mem_bus_if].rsp_valid;
								// Trace: src/VX_socket.sv:218:5
								assign l1_mem_arb_bus_if[0].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[0 + _mbase_mem_bus_if].rsp_data;
								// Trace: src/VX_socket.sv:219:5
								assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[0 + _mbase_mem_bus_if].rsp_ready = l1_mem_arb_bus_if[0].rsp_ready;
							end
							else begin : g_i
								// Trace: src/VX_socket.sv:221:13
								// expanded interface instance: l1_mem_arb_bus_if
								localparam _param_D5D25_DATA_SIZE = 64;
								localparam _param_D5D25_TAG_WIDTH = VX_gpu_pkg_L1_MEM_ARB_TAG_WIDTH;
								if (1) begin : l1_mem_arb_bus_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_bus_if.sv:2:15
									localparam DATA_SIZE = _param_D5D25_DATA_SIZE;
									// Trace: src/VX_mem_bus_if.sv:3:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:4:15
									localparam TAG_WIDTH = _param_D5D25_TAG_WIDTH;
									// Trace: src/VX_mem_bus_if.sv:5:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_mem_bus_if.sv:6:15
									localparam ADDR_WIDTH = 26;
									// Trace: src/VX_mem_bus_if.sv:8:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type tag_t
									// Trace: src/VX_mem_bus_if.sv:12:5
									// removed localparam type req_data_t
									// Trace: src/VX_mem_bus_if.sv:20:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_mem_bus_if.sv:24:5
									wire req_valid;
									// Trace: src/VX_mem_bus_if.sv:25:5
									wire [612:0] req_data;
									// Trace: src/VX_mem_bus_if.sv:26:5
									wire req_ready;
									// Trace: src/VX_mem_bus_if.sv:27:5
									wire rsp_valid;
									// Trace: src/VX_mem_bus_if.sv:28:5
									wire [518:0] rsp_data;
									// Trace: src/VX_mem_bus_if.sv:29:5
									wire rsp_ready;
									// Trace: src/VX_mem_bus_if.sv:30:5
									// Trace: src/VX_mem_bus_if.sv:38:5
								end
								// Trace: src/VX_socket.sv:226:5
								assign l1_mem_arb_bus_if.req_valid = dcache_mem_bus_if[i].req_valid;
								// Trace: src/VX_socket.sv:227:5
								assign l1_mem_arb_bus_if.req_data[612] = dcache_mem_bus_if[i].req_data[611];
								// Trace: src/VX_socket.sv:228:5
								assign l1_mem_arb_bus_if.req_data[611-:26] = dcache_mem_bus_if[i].req_data[610-:26];
								// Trace: src/VX_socket.sv:229:5
								assign l1_mem_arb_bus_if.req_data[585-:512] = dcache_mem_bus_if[i].req_data[584-:512];
								// Trace: src/VX_socket.sv:230:5
								assign l1_mem_arb_bus_if.req_data[73-:64] = dcache_mem_bus_if[i].req_data[72-:64];
								// Trace: src/VX_socket.sv:231:5
								assign l1_mem_arb_bus_if.req_data[9-:3] = dcache_mem_bus_if[i].req_data[8-:3];
								if (1) begin : genblk1
									if (1) begin : genblk1
										if (1) begin : genblk1
											// Trace: src/VX_socket.sv:235:17
											assign l1_mem_arb_bus_if.req_data[6-:7] = {dcache_mem_bus_if[i].req_data[5-:1], 1'b0, dcache_mem_bus_if[i].req_data[4-:5]};
										end
									end
								end
								// Trace: src/VX_socket.sv:249:5
								assign dcache_mem_bus_if[i].req_ready = l1_mem_arb_bus_if.req_ready;
								// Trace: src/VX_socket.sv:250:5
								assign dcache_mem_bus_if[i].rsp_valid = l1_mem_arb_bus_if.rsp_valid;
								// Trace: src/VX_socket.sv:251:5
								assign dcache_mem_bus_if[i].rsp_data[517-:512] = l1_mem_arb_bus_if.rsp_data[518-:512];
								if (1) begin : genblk2
									if (1) begin : genblk1
										if (1) begin : genblk1
											// Trace: src/VX_socket.sv:255:17
											assign dcache_mem_bus_if[i].rsp_data[5-:6] = {l1_mem_arb_bus_if.rsp_data[6-:1], l1_mem_arb_bus_if.rsp_data[4:0]};
										end
									end
								end
								// Trace: src/VX_socket.sv:269:5
								assign l1_mem_arb_bus_if.rsp_ready = dcache_mem_bus_if[i].rsp_ready;
								// Trace: src/VX_socket.sv:271:5
								assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_mem_bus_if].req_valid = l1_mem_arb_bus_if.req_valid;
								// Trace: src/VX_socket.sv:272:5
								assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_mem_bus_if].req_data = l1_mem_arb_bus_if.req_data;
								// Trace: src/VX_socket.sv:273:5
								assign l1_mem_arb_bus_if.req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_mem_bus_if].req_ready;
								// Trace: src/VX_socket.sv:274:5
								assign l1_mem_arb_bus_if.rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_mem_bus_if].rsp_valid;
								// Trace: src/VX_socket.sv:275:5
								assign l1_mem_arb_bus_if.rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_mem_bus_if].rsp_data;
								// Trace: src/VX_socket.sv:276:5
								assign Vortex.g_clusters[_gv_cluster_id_1].cluster.per_socket_mem_bus_if[i + _mbase_mem_bus_if].rsp_ready = l1_mem_arb_bus_if.rsp_ready;
							end
						end
						// Trace: src/VX_socket.sv:279:5
						wire [0:0] per_core_busy;
						// Trace: src/VX_socket.sv:280:5
						genvar _gv_core_id_1;
						localparam VX_gpu_pkg_VX_DCR_ADDR_WIDTH = 12;
						localparam VX_gpu_pkg_VX_DCR_DATA_WIDTH = 32;
						for (_gv_core_id_1 = 0; _gv_core_id_1 < 1; _gv_core_id_1 = _gv_core_id_1 + 1) begin : g_cores
							localparam core_id = _gv_core_id_1;
							// Trace: src/VX_socket.sv:281:5
							wire [0:0] core_reset;
							// Trace: src/VX_socket.sv:282:5
							VX_reset_relay #(
								.N(1),
								.MAX_FANOUT(0)
							) __core_reset(
								.clk(clk),
								.reset(reset),
								.reset_o(core_reset)
							);
							// Trace: src/VX_socket.sv:287:9
							// expanded interface instance: core_dcr_bus_if
							if (1) begin : core_dcr_bus_if
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_dcr_bus_if.sv:2:5
								wire write_valid;
								// Trace: src/VX_dcr_bus_if.sv:3:5
								localparam VX_gpu_pkg_VX_DCR_ADDR_WIDTH = 12;
								wire [11:0] write_addr;
								// Trace: src/VX_dcr_bus_if.sv:4:5
								localparam VX_gpu_pkg_VX_DCR_DATA_WIDTH = 32;
								wire [31:0] write_data;
								// Trace: src/VX_dcr_bus_if.sv:5:5
								// Trace: src/VX_dcr_bus_if.sv:10:5
							end
							if (1) begin : genblk1
								// Trace: src/VX_socket.sv:301:9
								assign {core_dcr_bus_if.write_valid, core_dcr_bus_if.write_addr, core_dcr_bus_if.write_data} = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket_dcr_bus_if.write_valid && 1'b1, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket_dcr_bus_if.write_addr, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket_dcr_bus_if.write_data};
							end
							// Trace: src/VX_socket.sv:304:9
							// expanded module instance: core
							localparam _bbase_588EE_dcache_bus_if = core_id * VX_gpu_pkg_DCACHE_NUM_REQS;
							localparam _bbase_588EE_icache_bus_if = core_id;
							localparam _param_588EE_CORE_ID = (SOCKET_ID * 1) + core_id;
							localparam _param_588EE_INSTANCE_ID = "";
							if (1) begin : core
								// removed import VX_gpu_pkg::*;
								// Trace: src/VX_core.sv:2:15
								localparam CORE_ID = _param_588EE_CORE_ID;
								// Trace: src/VX_core.sv:3:15
								localparam INSTANCE_ID = _param_588EE_INSTANCE_ID;
								// Trace: src/VX_core.sv:5:5
								wire clk;
								// Trace: src/VX_core.sv:6:5
								wire reset;
								// Trace: src/VX_core.sv:7:5
								// removed modport instance dcr_bus_if
								// Trace: src/VX_core.sv:8:5
								localparam VX_gpu_pkg_DCACHE_WORD_SIZE = 16;
								localparam VX_gpu_pkg_XLENB = 4;
								localparam VX_gpu_pkg_LSU_WORD_SIZE = VX_gpu_pkg_XLENB;
								localparam VX_gpu_pkg_DCACHE_CHANNELS = 1;
								localparam VX_gpu_pkg_DCACHE_NUM_REQS = 1;
								localparam _mbase_dcache_bus_if = _bbase_588EE_dcache_bus_if;
								// Trace: src/VX_core.sv:9:5
								localparam _mbase_icache_bus_if = _bbase_588EE_icache_bus_if;
								// Trace: src/VX_core.sv:10:5
								wire busy;
								// Trace: src/VX_core.sv:12:5
								// expanded interface instance: schedule_if
								if (1) begin : schedule_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_schedule_if.sv:2:5
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									localparam VX_gpu_pkg_PC_BITS = 30;
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type data_t
									// Trace: src/VX_schedule_if.sv:8:5
									wire valid;
									// Trace: src/VX_schedule_if.sv:9:5
									wire [36:0] data;
									// Trace: src/VX_schedule_if.sv:10:5
									wire ready;
									// Trace: src/VX_schedule_if.sv:11:5
									// Trace: src/VX_schedule_if.sv:16:5
								end
								// Trace: src/VX_core.sv:13:5
								// expanded interface instance: fetch_if
								if (1) begin : fetch_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_fetch_if.sv:2:5
									wire valid;
									// Trace: src/VX_fetch_if.sv:3:5
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									localparam VX_gpu_pkg_PC_BITS = 30;
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type VX_gpu_pkg_fetch_t
									wire [68:0] data;
									// Trace: src/VX_fetch_if.sv:4:5
									wire ready;
									// Trace: src/VX_fetch_if.sv:5:5
									// Trace: src/VX_fetch_if.sv:10:5
								end
								// Trace: src/VX_core.sv:14:5
								// expanded interface instance: decode_if
								if (1) begin : decode_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_decode_if.sv:2:5
									wire valid;
									// Trace: src/VX_decode_if.sv:3:5
									localparam VX_gpu_pkg_EX_SFU = 2;
									localparam VX_gpu_pkg_EX_FPU = 2;
									localparam VX_gpu_pkg_EX_TCU = 2;
									localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
									localparam VX_gpu_pkg_EX_BITS = 2;
									localparam VX_gpu_pkg_INST_OP_BITS = 4;
									localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									localparam VX_gpu_pkg_PC_BITS = 30;
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
									// removed localparam type VX_gpu_pkg_alu_args_t
									localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
									// removed localparam type VX_gpu_pkg_csr_args_t
									localparam VX_gpu_pkg_INST_FMT_BITS = 2;
									localparam VX_gpu_pkg_INST_FRM_BITS = 3;
									// removed localparam type VX_gpu_pkg_fpu_args_t
									localparam VX_gpu_pkg_OFFSET_BITS = 12;
									// removed localparam type VX_gpu_pkg_lsu_args_t
									// removed localparam type VX_gpu_pkg_wctl_args_t
									// removed localparam type VX_gpu_pkg_op_args_t
									localparam VX_gpu_pkg_REG_TYPES = 1;
									localparam VX_gpu_pkg_REG_TYPE_BITS = 1;
									localparam VX_gpu_pkg_RV_REGS_BITS = 5;
									// removed localparam type VX_gpu_pkg_reg_idx_t
									// removed localparam type VX_gpu_pkg_decode_t
									wire [107:0] data;
									// Trace: src/VX_decode_if.sv:4:5
									wire ready;
									// Trace: src/VX_decode_if.sv:5:5
									// Trace: src/VX_decode_if.sv:10:5
								end
								// Trace: src/VX_core.sv:15:5
								// expanded interface instance: sched_csr_if
								if (1) begin : sched_csr_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_sched_csr_if.sv:2:5
									localparam VX_gpu_pkg_PERF_CTR_BITS = 44;
									wire [43:0] cycles;
									// Trace: src/VX_sched_csr_if.sv:3:5
									wire [3:0] active_warps;
									// Trace: src/VX_sched_csr_if.sv:4:5
									wire [15:0] thread_masks;
									// Trace: src/VX_sched_csr_if.sv:5:5
									wire alm_empty;
									// Trace: src/VX_sched_csr_if.sv:6:5
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									wire [1:0] alm_empty_wid;
									// Trace: src/VX_sched_csr_if.sv:7:5
									wire unlock_warp;
									// Trace: src/VX_sched_csr_if.sv:8:5
									wire [1:0] unlock_wid;
									// Trace: src/VX_sched_csr_if.sv:9:5
									// Trace: src/VX_sched_csr_if.sv:18:5
								end
								// Trace: src/VX_core.sv:16:5
								// expanded interface instance: decode_sched_if
								if (1) begin : decode_sched_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_decode_sched_if.sv:2:5
									wire valid;
									// Trace: src/VX_decode_sched_if.sv:3:5
									wire unlock;
									// Trace: src/VX_decode_sched_if.sv:4:5
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									wire [1:0] wid;
									// Trace: src/VX_decode_sched_if.sv:5:5
									// Trace: src/VX_decode_sched_if.sv:10:5
								end
								// Trace: src/VX_core.sv:17:5
								// expanded interface instance: issue_sched_if
								genvar _arr_E332A;
								for (_arr_E332A = 0; _arr_E332A <= 0; _arr_E332A = _arr_E332A + 1) begin : issue_sched_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_issue_sched_if.sv:2:5
									localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
									localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
									localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
									wire [1:0] wis;
									// Trace: src/VX_issue_sched_if.sv:3:5
									wire valid;
									// Trace: src/VX_issue_sched_if.sv:4:5
									// Trace: src/VX_issue_sched_if.sv:8:5
								end
								// Trace: src/VX_core.sv:18:5
								// expanded interface instance: commit_sched_if
								if (1) begin : commit_sched_if
									// Trace: src/VX_commit_sched_if.sv:2:5
									wire [3:0] committed_warps;
									// Trace: src/VX_commit_sched_if.sv:3:5
									// Trace: src/VX_commit_sched_if.sv:6:5
								end
								// Trace: src/VX_core.sv:19:5
								// expanded interface instance: commit_csr_if
								if (1) begin : commit_csr_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_commit_csr_if.sv:2:5
									localparam VX_gpu_pkg_PERF_CTR_BITS = 44;
									wire [43:0] instret;
									// Trace: src/VX_commit_csr_if.sv:3:5
									// Trace: src/VX_commit_csr_if.sv:6:5
								end
								// Trace: src/VX_core.sv:20:5
								// expanded interface instance: branch_ctl_if
								genvar _arr_DDFE6;
								for (_arr_DDFE6 = 0; _arr_DDFE6 <= 0; _arr_DDFE6 = _arr_DDFE6 + 1) begin : branch_ctl_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_branch_ctl_if.sv:2:5
									wire valid;
									// Trace: src/VX_branch_ctl_if.sv:3:5
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									wire [1:0] wid;
									// Trace: src/VX_branch_ctl_if.sv:4:5
									wire taken;
									// Trace: src/VX_branch_ctl_if.sv:5:5
									localparam VX_gpu_pkg_PC_BITS = 30;
									wire [29:0] dest;
									// Trace: src/VX_branch_ctl_if.sv:6:5
									// Trace: src/VX_branch_ctl_if.sv:12:5
								end
								// Trace: src/VX_core.sv:21:5
								// expanded interface instance: warp_ctl_if
								if (1) begin : warp_ctl_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_warp_ctl_if.sv:2:5
									wire valid;
									// Trace: src/VX_warp_ctl_if.sv:3:5
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									wire [1:0] wid;
									// Trace: src/VX_warp_ctl_if.sv:4:5
									// removed localparam type VX_gpu_pkg_tmc_t
									wire [4:0] tmc;
									// Trace: src/VX_warp_ctl_if.sv:5:5
									localparam VX_gpu_pkg_PC_BITS = 30;
									// removed localparam type VX_gpu_pkg_wspawn_t
									wire [34:0] wspawn;
									// Trace: src/VX_warp_ctl_if.sv:6:5
									// removed localparam type VX_gpu_pkg_split_t
									wire [39:0] split;
									// Trace: src/VX_warp_ctl_if.sv:7:5
									localparam VX_gpu_pkg_DV_STACK_SIZE = 3;
									localparam VX_gpu_pkg_DV_STACK_SIZEW = 2;
									// removed localparam type VX_gpu_pkg_join_t
									wire [2:0] sjoin;
									// Trace: src/VX_warp_ctl_if.sv:8:5
									localparam VX_gpu_pkg_NB_BITS = 1;
									localparam VX_gpu_pkg_NB_WIDTH = VX_gpu_pkg_NB_BITS;
									// removed localparam type VX_gpu_pkg_barrier_t
									wire [5:0] barrier;
									// Trace: src/VX_warp_ctl_if.sv:9:5
									wire [1:0] dvstack_wid;
									// Trace: src/VX_warp_ctl_if.sv:10:5
									wire [1:0] dvstack_ptr;
									// Trace: src/VX_warp_ctl_if.sv:11:5
									// Trace: src/VX_warp_ctl_if.sv:22:5
								end
								// Trace: src/VX_core.sv:22:5
								localparam VX_gpu_pkg_EX_SFU = 2;
								localparam VX_gpu_pkg_EX_FPU = 2;
								localparam VX_gpu_pkg_EX_TCU = 2;
								localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
								// expanded interface instance: dispatch_if
								genvar _arr_B1D72;
								for (_arr_B1D72 = 0; _arr_B1D72 <= 2; _arr_B1D72 = _arr_B1D72 + 1) begin : dispatch_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_dispatch_if.sv:2:5
									wire valid;
									// Trace: src/VX_dispatch_if.sv:3:5
									localparam VX_gpu_pkg_INST_ALU_BITS = 4;
									localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
									localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
									localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
									localparam VX_gpu_pkg_REG_TYPES = 1;
									localparam VX_gpu_pkg_RV_REGS = 32;
									localparam VX_gpu_pkg_NUM_REGS = 32;
									localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
									localparam VX_gpu_pkg_PC_BITS = 30;
									localparam VX_gpu_pkg_SIMD_COUNT = 1;
									localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
									localparam VX_gpu_pkg_SIMD_IDX_W = 1;
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
									// removed localparam type VX_gpu_pkg_alu_args_t
									localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
									// removed localparam type VX_gpu_pkg_csr_args_t
									localparam VX_gpu_pkg_INST_FMT_BITS = 2;
									localparam VX_gpu_pkg_INST_FRM_BITS = 3;
									// removed localparam type VX_gpu_pkg_fpu_args_t
									localparam VX_gpu_pkg_OFFSET_BITS = 12;
									// removed localparam type VX_gpu_pkg_lsu_args_t
									// removed localparam type VX_gpu_pkg_wctl_args_t
									// removed localparam type VX_gpu_pkg_op_args_t
									// removed localparam type VX_gpu_pkg_dispatch_t
									wire [470:0] data;
									// Trace: src/VX_dispatch_if.sv:4:5
									wire ready;
									// Trace: src/VX_dispatch_if.sv:5:5
									// Trace: src/VX_dispatch_if.sv:10:5
								end
								// Trace: src/VX_core.sv:23:5
								// expanded interface instance: commit_if
								genvar _arr_56FA2;
								for (_arr_56FA2 = 0; _arr_56FA2 <= 2; _arr_56FA2 = _arr_56FA2 + 1) begin : commit_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_commit_if.sv:2:5
									wire valid;
									// Trace: src/VX_commit_if.sv:3:5
									localparam VX_gpu_pkg_REG_TYPES = 1;
									localparam VX_gpu_pkg_RV_REGS = 32;
									localparam VX_gpu_pkg_NUM_REGS = 32;
									localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									localparam VX_gpu_pkg_PC_BITS = 30;
									localparam VX_gpu_pkg_SIMD_COUNT = 1;
									localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
									localparam VX_gpu_pkg_SIMD_IDX_W = 1;
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type VX_gpu_pkg_commit_t
									wire [173:0] data;
									// Trace: src/VX_commit_if.sv:4:5
									wire ready;
									// Trace: src/VX_commit_if.sv:5:5
									// Trace: src/VX_commit_if.sv:10:5
								end
								// Trace: src/VX_core.sv:24:5
								// expanded interface instance: writeback_if
								genvar _arr_8BCF0;
								for (_arr_8BCF0 = 0; _arr_8BCF0 <= 0; _arr_8BCF0 = _arr_8BCF0 + 1) begin : writeback_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_writeback_if.sv:2:5
									wire valid;
									// Trace: src/VX_writeback_if.sv:3:5
									localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
									localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
									localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
									localparam VX_gpu_pkg_REG_TYPES = 1;
									localparam VX_gpu_pkg_RV_REGS = 32;
									localparam VX_gpu_pkg_NUM_REGS = 32;
									localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
									localparam VX_gpu_pkg_PC_BITS = 30;
									localparam VX_gpu_pkg_SIMD_COUNT = 1;
									localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
									localparam VX_gpu_pkg_SIMD_IDX_W = 1;
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type VX_gpu_pkg_writeback_t
									wire [172:0] data;
									// Trace: src/VX_writeback_if.sv:4:5
									// Trace: src/VX_writeback_if.sv:8:5
								end
								// Trace: src/VX_core.sv:25:5
								localparam VX_gpu_pkg_LSU_MEM_BATCHES = 1;
								localparam VX_gpu_pkg_LSU_TAG_ID_BITS = 1;
								localparam VX_gpu_pkg_UUID_WIDTH = 1;
								localparam VX_gpu_pkg_LSU_TAG_WIDTH = 2;
								// expanded interface instance: lsu_mem_if
								localparam _param_DD8FC_NUM_LANES = 4;
								localparam _param_DD8FC_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
								localparam _param_DD8FC_TAG_WIDTH = VX_gpu_pkg_LSU_TAG_WIDTH;
								genvar _arr_DD8FC;
								for (_arr_DD8FC = 0; _arr_DD8FC <= 0; _arr_DD8FC = _arr_DD8FC + 1) begin : lsu_mem_if
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_lsu_mem_if.sv:2:15
									localparam NUM_LANES = _param_DD8FC_NUM_LANES;
									// Trace: src/VX_lsu_mem_if.sv:3:15
									localparam DATA_SIZE = _param_DD8FC_DATA_SIZE;
									// Trace: src/VX_lsu_mem_if.sv:4:15
									localparam TAG_WIDTH = _param_DD8FC_TAG_WIDTH;
									// Trace: src/VX_lsu_mem_if.sv:5:15
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
									// Trace: src/VX_lsu_mem_if.sv:6:15
									localparam MEM_ADDR_WIDTH = 32;
									// Trace: src/VX_lsu_mem_if.sv:7:15
									localparam ADDR_WIDTH = 30;
									// Trace: src/VX_lsu_mem_if.sv:9:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type tag_t
									// Trace: src/VX_lsu_mem_if.sv:13:5
									// removed localparam type req_data_t
									// Trace: src/VX_lsu_mem_if.sv:22:5
									// removed localparam type rsp_data_t
									// Trace: src/VX_lsu_mem_if.sv:27:5
									wire req_valid;
									// Trace: src/VX_lsu_mem_if.sv:28:5
									wire [282:0] req_data;
									// Trace: src/VX_lsu_mem_if.sv:29:5
									wire req_ready;
									// Trace: src/VX_lsu_mem_if.sv:30:5
									wire rsp_valid;
									// Trace: src/VX_lsu_mem_if.sv:31:5
									wire [133:0] rsp_data;
									// Trace: src/VX_lsu_mem_if.sv:32:5
									wire rsp_ready;
									// Trace: src/VX_lsu_mem_if.sv:33:5
									// Trace: src/VX_lsu_mem_if.sv:41:5
								end
								// Trace: src/VX_core.sv:30:5
								// removed localparam type VX_gpu_pkg_base_dcrs_t
								wire [71:0] base_dcrs;
								// Trace: src/VX_core.sv:31:5
								// expanded module instance: dcr_data
								if (1) begin : dcr_data
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_dcr_data.sv:2:5
									wire clk;
									// Trace: src/VX_dcr_data.sv:3:5
									wire reset;
									// Trace: src/VX_dcr_data.sv:4:5
									// removed modport instance dcr_bus_if
									// Trace: src/VX_dcr_data.sv:5:5
									// removed localparam type VX_gpu_pkg_base_dcrs_t
									wire [71:0] base_dcrs;
									// Trace: src/VX_dcr_data.sv:7:5
									reg [71:0] dcrs;
									// Trace: src/VX_dcr_data.sv:8:5
									always @(posedge clk)
										// Trace: src/VX_dcr_data.sv:9:8
										if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core_dcr_bus_if.write_valid)
											// Trace: src/VX_dcr_data.sv:10:13
											case (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core_dcr_bus_if.write_addr)
												12'h001:
													// Trace: src/VX_dcr_data.sv:11:23
													dcrs[71:40] <= Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core_dcr_bus_if.write_data;
												12'h003:
													// Trace: src/VX_dcr_data.sv:12:23
													dcrs[39:8] <= Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core_dcr_bus_if.write_data;
												12'h005:
													// Trace: src/VX_dcr_data.sv:13:23
													dcrs[7-:8] <= Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core_dcr_bus_if.write_data[7:0];
												default:
													;
											endcase
									// Trace: src/VX_dcr_data.sv:18:5
									assign base_dcrs = dcrs;
								end
								assign dcr_data.clk = clk;
								assign dcr_data.reset = reset;
								assign base_dcrs = dcr_data.base_dcrs;
								// Trace: src/VX_core.sv:38:5
								// expanded module instance: schedule
								localparam _bbase_45092_branch_ctl_if = 0;
								localparam _bbase_45092_issue_sched_if = 0;
								localparam _param_45092_INSTANCE_ID = "";
								localparam _param_45092_CORE_ID = CORE_ID;
								if (1) begin : schedule
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_schedule.sv:2:15
									localparam INSTANCE_ID = _param_45092_INSTANCE_ID;
									// Trace: src/VX_schedule.sv:3:15
									localparam CORE_ID = _param_45092_CORE_ID;
									// Trace: src/VX_schedule.sv:5:5
									wire clk;
									// Trace: src/VX_schedule.sv:6:5
									wire reset;
									// Trace: src/VX_schedule.sv:7:5
									// removed localparam type VX_gpu_pkg_base_dcrs_t
									wire [71:0] base_dcrs;
									// Trace: src/VX_schedule.sv:8:5
									// removed modport instance warp_ctl_if
									// Trace: src/VX_schedule.sv:9:5
									localparam _mbase_branch_ctl_if = 0;
									// Trace: src/VX_schedule.sv:10:5
									// removed modport instance decode_sched_if
									// Trace: src/VX_schedule.sv:11:5
									localparam _mbase_issue_sched_if = 0;
									// Trace: src/VX_schedule.sv:12:5
									// removed modport instance commit_sched_if
									// Trace: src/VX_schedule.sv:13:5
									// removed modport instance schedule_if
									// Trace: src/VX_schedule.sv:14:5
									// removed modport instance sched_csr_if
									// Trace: src/VX_schedule.sv:15:5
									wire busy;
									// Trace: src/VX_schedule.sv:17:5
									reg [3:0] active_warps;
									reg [3:0] active_warps_n;
									// Trace: src/VX_schedule.sv:18:5
									reg [3:0] stalled_warps;
									reg [3:0] stalled_warps_n;
									// Trace: src/VX_schedule.sv:19:5
									reg [15:0] thread_masks;
									reg [15:0] thread_masks_n;
									// Trace: src/VX_schedule.sv:20:5
									localparam VX_gpu_pkg_PC_BITS = 30;
									reg [119:0] warp_pcs;
									reg [119:0] warp_pcs_n;
									// Trace: src/VX_schedule.sv:21:5
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									wire [1:0] schedule_wid;
									// Trace: src/VX_schedule.sv:22:5
									wire [3:0] schedule_tmask;
									// Trace: src/VX_schedule.sv:23:5
									wire [29:0] schedule_pc;
									// Trace: src/VX_schedule.sv:24:5
									wire schedule_valid;
									// Trace: src/VX_schedule.sv:25:5
									wire schedule_ready;
									// Trace: src/VX_schedule.sv:26:5
									wire join_valid;
									// Trace: src/VX_schedule.sv:27:5
									wire join_is_dvg;
									// Trace: src/VX_schedule.sv:28:5
									wire join_is_else;
									// Trace: src/VX_schedule.sv:29:5
									wire [1:0] join_wid;
									// Trace: src/VX_schedule.sv:30:5
									wire [3:0] join_tmask;
									// Trace: src/VX_schedule.sv:31:5
									wire [29:0] join_pc;
									// Trace: src/VX_schedule.sv:32:5
									localparam VX_gpu_pkg_PERF_CTR_BITS = 44;
									reg [43:0] cycles;
									// Trace: src/VX_schedule.sv:33:5
									wire schedule_fire = schedule_valid && schedule_ready;
									// Trace: src/VX_schedule.sv:34:5
									wire schedule_if_fire = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.ready;
									// Trace: src/VX_schedule.sv:35:5
									wire [0:0] branch_valid;
									// Trace: src/VX_schedule.sv:36:5
									wire [1:0] branch_wid;
									// Trace: src/VX_schedule.sv:37:5
									wire [0:0] branch_taken;
									// Trace: src/VX_schedule.sv:38:5
									wire [29:0] branch_dest;
									// Trace: src/VX_schedule.sv:39:5
									genvar _gv_i_5;
									for (_gv_i_5 = 0; _gv_i_5 < 1; _gv_i_5 = _gv_i_5 + 1) begin : g_branch_init
										localparam i = _gv_i_5;
										// Trace: src/VX_schedule.sv:40:9
										assign branch_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[i + _mbase_branch_ctl_if].valid;
										// Trace: src/VX_schedule.sv:41:9
										assign branch_wid[i * 2+:2] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[i + _mbase_branch_ctl_if].wid;
										// Trace: src/VX_schedule.sv:42:9
										assign branch_taken[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[i + _mbase_branch_ctl_if].taken;
										// Trace: src/VX_schedule.sv:43:9
										assign branch_dest[i * 30+:30] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[i + _mbase_branch_ctl_if].dest;
									end
									// Trace: src/VX_schedule.sv:45:5
									reg [7:0] barrier_masks;
									reg [7:0] barrier_masks_n;
									// Trace: src/VX_schedule.sv:46:5
									reg [3:0] barrier_ctrs;
									reg [3:0] barrier_ctrs_n;
									// Trace: src/VX_schedule.sv:47:5
									reg [3:0] barrier_stalls;
									reg [3:0] barrier_stalls_n;
									// Trace: src/VX_schedule.sv:48:5
									reg [3:0] curr_barrier_mask_p1;
									// Trace: src/VX_schedule.sv:49:5
									// removed localparam type VX_gpu_pkg_wspawn_t
									reg [34:0] wspawn;
									// Trace: src/VX_schedule.sv:50:5
									reg [1:0] wspawn_wid;
									// Trace: src/VX_schedule.sv:51:5
									reg is_single_warp;
									// Trace: src/VX_schedule.sv:52:5
									wire [2:0] active_warps_cnt;
									// Trace: src/VX_schedule.sv:53:5
									VX_popcount #(
										.N(4),
										.MODEL(1)
									) __pop_count_ex104(
										.data_in(active_warps),
										.data_out(active_warps_cnt)
									);
									// Trace: src/VX_schedule.sv:60:5
									function automatic [29:0] VX_gpu_pkg_from_fullPC;
										// Trace: src/VX_gpu_pkg.sv:30:56
										input reg [31:0] pc;
										// Trace: src/VX_gpu_pkg.sv:31:9
										VX_gpu_pkg_from_fullPC = sv2v_cast_30(pc >> 2);
									endfunction
									always @(*) begin
										// Trace: src/VX_schedule.sv:61:9
										active_warps_n = active_warps;
										// Trace: src/VX_schedule.sv:62:9
										stalled_warps_n = stalled_warps;
										// Trace: src/VX_schedule.sv:63:9
										thread_masks_n = thread_masks;
										// Trace: src/VX_schedule.sv:64:9
										barrier_masks_n = barrier_masks;
										// Trace: src/VX_schedule.sv:65:9
										barrier_ctrs_n = barrier_ctrs;
										// Trace: src/VX_schedule.sv:66:9
										barrier_stalls_n = barrier_stalls;
										// Trace: src/VX_schedule.sv:67:9
										warp_pcs_n = warp_pcs;
										// Trace: src/VX_schedule.sv:68:9
										if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.unlock)
											// Trace: src/VX_schedule.sv:69:13
											stalled_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.wid] = 0;
										if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.unlock_warp)
											// Trace: src/VX_schedule.sv:72:13
											stalled_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.unlock_wid] = 0;
										if (wspawn[34] && is_single_warp) begin
											// Trace: src/VX_schedule.sv:75:13
											active_warps_n = active_warps_n | wspawn[33-:4];
											// Trace: src/VX_schedule.sv:76:13
											begin : sv2v_autoblock_3
												// Trace: src/VX_schedule.sv:76:18
												integer i;
												// Trace: src/VX_schedule.sv:76:18
												for (i = 0; i < 4; i = i + 1)
													begin
														// Trace: src/VX_schedule.sv:77:17
														if (wspawn[30 + i]) begin
															// Trace: src/VX_schedule.sv:78:21
															thread_masks_n[i * 4] = 1;
															// Trace: src/VX_schedule.sv:79:21
															warp_pcs_n[i * 30+:30] = wspawn[29-:30];
														end
													end
											end
											// Trace: src/VX_schedule.sv:82:13
											stalled_warps_n[wspawn_wid] = 0;
										end
										if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.tmc[4]) begin
											// Trace: src/VX_schedule.sv:85:13
											active_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.tmc[3-:4] != 0;
											// Trace: src/VX_schedule.sv:86:13
											thread_masks_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid * 4+:4] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.tmc[3-:4];
											// Trace: src/VX_schedule.sv:87:13
											stalled_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid] = 0;
										end
										if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.split[39]) begin
											// Trace: src/VX_schedule.sv:90:13
											if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.split[38])
												// Trace: src/VX_schedule.sv:91:17
												thread_masks_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid * 4+:4] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.split[37-:4];
											// Trace: src/VX_schedule.sv:93:13
											stalled_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid] = 0;
										end
										if (join_valid) begin
											// Trace: src/VX_schedule.sv:96:13
											if (join_is_dvg) begin
												// Trace: src/VX_schedule.sv:97:17
												if (join_is_else)
													// Trace: src/VX_schedule.sv:98:21
													warp_pcs_n[join_wid * 30+:30] = join_pc;
												// Trace: src/VX_schedule.sv:100:17
												thread_masks_n[join_wid * 4+:4] = join_tmask;
											end
											// Trace: src/VX_schedule.sv:102:13
											stalled_warps_n[join_wid] = 0;
										end
										// Trace: src/VX_schedule.sv:104:9
										curr_barrier_mask_p1 = barrier_masks[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 4+:4];
										// Trace: src/VX_schedule.sv:105:9
										curr_barrier_mask_p1[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid] = 1;
										if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[5]) begin
											begin
												// Trace: src/VX_schedule.sv:107:13
												if (~Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[0]) begin
													begin
														// Trace: src/VX_schedule.sv:108:17
														if (~Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[3] && (barrier_ctrs[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 2+:2] == sv2v_cast_2(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[2-:2]))) begin
															// Trace: src/VX_schedule.sv:110:21
															barrier_ctrs_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 2+:2] = 1'sb0;
															// Trace: src/VX_schedule.sv:111:21
															barrier_masks_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 4+:4] = 1'sb0;
															// Trace: src/VX_schedule.sv:112:21
															stalled_warps_n = stalled_warps_n & ~barrier_masks[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 4+:4];
															// Trace: src/VX_schedule.sv:113:21
															stalled_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid] = 0;
														end
														else begin
															// Trace: src/VX_schedule.sv:115:21
															barrier_ctrs_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 2+:2] = barrier_ctrs[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 2+:2] + 2'sd1;
															// Trace: src/VX_schedule.sv:116:21
															barrier_masks_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier[4-:1] * 4+:4] = curr_barrier_mask_p1;
														end
													end
												end
												else
													// Trace: src/VX_schedule.sv:119:17
													stalled_warps_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid] = 0;
											end
										end
										begin : sv2v_autoblock_4
											// Trace: src/VX_schedule.sv:122:14
											integer i;
											// Trace: src/VX_schedule.sv:122:14
											for (i = 0; i < 1; i = i + 1)
												begin
													// Trace: src/VX_schedule.sv:123:13
													if (branch_valid[i]) begin
														// Trace: src/VX_schedule.sv:124:17
														if (branch_taken[i])
															// Trace: src/VX_schedule.sv:125:21
															warp_pcs_n[branch_wid[i * 2+:2] * 30+:30] = branch_dest[i * 30+:30];
														// Trace: src/VX_schedule.sv:127:17
														stalled_warps_n[branch_wid[i * 2+:2]] = 0;
													end
												end
										end
										if (schedule_fire)
											// Trace: src/VX_schedule.sv:131:13
											stalled_warps_n[schedule_wid] = 1;
										if (schedule_if_fire)
											// Trace: src/VX_schedule.sv:134:13
											warp_pcs_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[35-:2] * 30+:30] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[29-:30] + VX_gpu_pkg_from_fullPC(32'sd4);
									end
									// Trace: src/VX_schedule.sv:137:5
									always @(posedge clk)
										// Trace: src/VX_schedule.sv:138:9
										if (reset) begin
											// Trace: src/VX_schedule.sv:139:13
											barrier_masks <= 1'sb0;
											// Trace: src/VX_schedule.sv:140:13
											barrier_ctrs <= 1'sb0;
											// Trace: src/VX_schedule.sv:141:13
											stalled_warps <= 1'sb0;
											// Trace: src/VX_schedule.sv:142:13
											warp_pcs <= 1'sb0;
											// Trace: src/VX_schedule.sv:143:13
											active_warps <= 1'sb0;
											// Trace: src/VX_schedule.sv:144:13
											thread_masks <= 1'sb0;
											// Trace: src/VX_schedule.sv:145:13
											barrier_stalls <= 1'sb0;
											// Trace: src/VX_schedule.sv:146:13
											cycles <= 1'sb0;
											// Trace: src/VX_schedule.sv:147:13
											wspawn[34] <= 0;
											// Trace: src/VX_schedule.sv:148:13
											warp_pcs[0+:30] <= VX_gpu_pkg_from_fullPC(base_dcrs[71-:32]);
											// Trace: src/VX_schedule.sv:149:13
											active_warps[0] <= 1;
											// Trace: src/VX_schedule.sv:150:13
											thread_masks[0] <= 1;
											// Trace: src/VX_schedule.sv:151:13
											is_single_warp <= 1;
										end
										else begin
											// Trace: src/VX_schedule.sv:153:13
											active_warps <= active_warps_n;
											// Trace: src/VX_schedule.sv:154:13
											stalled_warps <= stalled_warps_n;
											// Trace: src/VX_schedule.sv:155:13
											thread_masks <= thread_masks_n;
											// Trace: src/VX_schedule.sv:156:13
											warp_pcs <= warp_pcs_n;
											// Trace: src/VX_schedule.sv:157:13
											barrier_masks <= barrier_masks_n;
											// Trace: src/VX_schedule.sv:158:13
											barrier_ctrs <= barrier_ctrs_n;
											// Trace: src/VX_schedule.sv:159:13
											barrier_stalls <= barrier_stalls_n;
											// Trace: src/VX_schedule.sv:160:13
											is_single_warp <= active_warps_cnt == sv2v_cast_22555_signed(1);
											// Trace: src/VX_schedule.sv:161:13
											if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wspawn[34]) begin
												// Trace: src/VX_schedule.sv:162:17
												wspawn[34] <= 1;
												// Trace: src/VX_schedule.sv:163:17
												wspawn[33-:4] <= Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wspawn[33-:4];
												// Trace: src/VX_schedule.sv:164:17
												wspawn[29-:30] <= Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wspawn[29-:30];
												// Trace: src/VX_schedule.sv:165:17
												wspawn_wid <= Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid;
											end
											if (wspawn[34] && is_single_warp)
												// Trace: src/VX_schedule.sv:168:17
												wspawn[34] <= 0;
											if (busy)
												// Trace: src/VX_schedule.sv:171:17
												cycles <= cycles + 1;
										end
									// Trace: src/VX_schedule.sv:175:5
									VX_split_join #(
										.INSTANCE_ID(""),
										.OUT_REG(1)
									) split_join(
										.clk(clk),
										.reset(reset),
										.valid(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.valid),
										.wid(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid),
										.split(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.split),
										.sjoin(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.sjoin),
										.join_valid(join_valid),
										.join_is_dvg(join_is_dvg),
										.join_is_else(join_is_else),
										.join_wid(join_wid),
										.join_tmask(join_tmask),
										.join_pc(join_pc),
										.stack_wid(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.dvstack_wid),
										.stack_ptr(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.dvstack_ptr)
									);
									// Trace: src/VX_schedule.sv:194:5
									wire [3:0] ready_warps = active_warps & ~stalled_warps;
									// Trace: src/VX_schedule.sv:195:5
									VX_priority_encoder #(.N(4)) wid_select(
										.data_in(ready_warps),
										.index_out(schedule_wid),
										.valid_out(schedule_valid),
										.onehot_out()
									);
									// Trace: src/VX_schedule.sv:203:5
									wire [135:0] schedule_data;
									// Trace: src/VX_schedule.sv:204:5
									genvar _gv_i_6;
									for (_gv_i_6 = 0; _gv_i_6 < 4; _gv_i_6 = _gv_i_6 + 1) begin : g_schedule_data
										localparam i = _gv_i_6;
										// Trace: src/VX_schedule.sv:205:9
										assign schedule_data[i * 34+:34] = {thread_masks[i * 4+:4], warp_pcs[i * 30+:30]};
									end
									// Trace: src/VX_schedule.sv:207:5
									assign {schedule_tmask, schedule_pc} = {schedule_data[(schedule_wid * 34) + 33-:4], schedule_data[(schedule_wid * 34) + 29-:30]};
									// Trace: src/VX_schedule.sv:211:5
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									wire [0:0] instr_uuid;
									// Trace: src/VX_schedule.sv:212:5
									assign instr_uuid = 1'sb0;
									// Trace: src/VX_schedule.sv:213:5
									VX_elastic_buffer #(
										.DATAW(37),
										.SIZE(2),
										.OUT_REG(1)
									) out_buf(
										.clk(clk),
										.reset(reset),
										.valid_in(schedule_valid),
										.ready_in(schedule_ready),
										.data_in({schedule_tmask, schedule_pc, schedule_wid, instr_uuid}),
										.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[33-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[29-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[35-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[36-:1]}),
										.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.valid),
										.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.ready)
									);
									// Trace: src/VX_schedule.sv:227:5
									wire [3:0] pending_warp_empty;
									// Trace: src/VX_schedule.sv:228:5
									wire [3:0] pending_warp_alm_empty;
									// Trace: src/VX_schedule.sv:229:5
									genvar _gv_i_7;
									localparam VX_gpu_pkg_ISSUE_ISW_BITS = 0;
									localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
									function automatic [0:0] VX_gpu_pkg_wid_to_isw;
										// Trace: src/VX_gpu_pkg.sv:276:9
										input reg [1:0] wid;
										// Trace: src/VX_gpu_pkg.sv:278:9
										begin
											// Trace: src/VX_gpu_pkg.sv:281:13
											VX_gpu_pkg_wid_to_isw = 0;
										end
									endfunction
									localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
									localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
									localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
									function automatic [1:0] VX_gpu_pkg_wid_to_wis;
										// Trace: src/VX_gpu_pkg.sv:285:9
										input reg [1:0] wid;
										// Trace: src/VX_gpu_pkg.sv:287:9
										begin
											// Trace: src/VX_gpu_pkg.sv:288:13
											VX_gpu_pkg_wid_to_wis = wid >> VX_gpu_pkg_ISSUE_ISW_BITS;
										end
									endfunction
									for (_gv_i_7 = 0; _gv_i_7 < 4; _gv_i_7 = _gv_i_7 + 1) begin : g_pending_sizes
										localparam i = _gv_i_7;
										// Trace: src/VX_schedule.sv:230:9
										localparam isw = VX_gpu_pkg_wid_to_isw(i);
										// Trace: src/VX_schedule.sv:231:9
										localparam wis = VX_gpu_pkg_wid_to_wis(i);
										// Trace: src/VX_schedule.sv:232:9
										VX_pending_size #(
											.SIZE(4096),
											.ALM_EMPTY(1)
										) counter(
											.clk(clk),
											.reset(reset),
											.incr(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue_sched_if[isw + _mbase_issue_sched_if].valid && (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue_sched_if[isw + _mbase_issue_sched_if].wis == wis)),
											.decr(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_sched_if.committed_warps[i]),
											.empty(pending_warp_empty[i]),
											.alm_empty(pending_warp_alm_empty[i]),
											.full(),
											.alm_full(),
											.size()
										);
									end
									// Trace: src/VX_schedule.sv:247:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.alm_empty = pending_warp_alm_empty[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.alm_empty_wid];
									// Trace: src/VX_schedule.sv:248:5
									wire no_pending_instr = &pending_warp_empty;
									// Trace: src/VX_schedule.sv:249:5
									VX_pipe_register #(
										.DATAW(1),
										.RESETW(1),
										.DEPTH(1)
									) __buffer_ex390(
										.clk(clk),
										.reset(reset),
										.enable(1'b1),
										.data_in((active_warps != 0) || ~no_pending_instr),
										.data_out(busy)
									);
									// Trace: src/VX_schedule.sv:260:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.cycles = cycles;
									// Trace: src/VX_schedule.sv:261:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.active_warps = active_warps;
									// Trace: src/VX_schedule.sv:262:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.thread_masks = thread_masks;
									// Trace: src/VX_schedule.sv:263:5
									reg [31:0] timeout_ctr;
									// Trace: src/VX_schedule.sv:264:5
									reg timeout_enable;
									// Trace: src/VX_schedule.sv:265:5
									always @(posedge clk)
										// Trace: src/VX_schedule.sv:266:9
										if (reset) begin
											// Trace: src/VX_schedule.sv:267:13
											timeout_ctr <= 1'sb0;
											// Trace: src/VX_schedule.sv:268:13
											timeout_enable <= 0;
										end
										else begin
											// Trace: src/VX_schedule.sv:270:13
											if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.unlock)
												// Trace: src/VX_schedule.sv:271:17
												timeout_enable <= 1;
											if ((timeout_enable && (active_warps != 0)) && (active_warps == stalled_warps))
												// Trace: src/VX_schedule.sv:274:17
												timeout_ctr <= timeout_ctr + 1;
											else if ((active_warps == 0) || (active_warps != stalled_warps))
												// Trace: src/VX_schedule.sv:276:17
												timeout_ctr <= 1'sb0;
										end
								end
								assign schedule.clk = clk;
								assign schedule.reset = reset;
								assign schedule.base_dcrs = base_dcrs;
								assign busy = schedule.busy;
								// Trace: src/VX_core.sv:54:5
								// expanded module instance: fetch
								localparam _bbase_852F6_icache_bus_if = core_id;
								localparam _param_852F6_INSTANCE_ID = "";
								if (1) begin : fetch
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_fetch.sv:2:15
									localparam INSTANCE_ID = _param_852F6_INSTANCE_ID;
									// Trace: src/VX_fetch.sv:4:5
									wire clk;
									// Trace: src/VX_fetch.sv:5:5
									wire reset;
									// Trace: src/VX_fetch.sv:6:5
									localparam _mbase_icache_bus_if = _bbase_852F6_icache_bus_if;
									// Trace: src/VX_fetch.sv:7:5
									// removed modport instance schedule_if
									// Trace: src/VX_fetch.sv:8:5
									// removed modport instance fetch_if
									// Trace: src/VX_fetch.sv:10:5
									wire icache_req_valid;
									// Trace: src/VX_fetch.sv:11:5
									localparam VX_gpu_pkg_ICACHE_WORD_SIZE = 4;
									localparam VX_gpu_pkg_ICACHE_ADDR_WIDTH = 30;
									wire [29:0] icache_req_addr;
									// Trace: src/VX_fetch.sv:12:5
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									localparam VX_gpu_pkg_ICACHE_TAG_ID_BITS = VX_gpu_pkg_NW_WIDTH;
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									localparam VX_gpu_pkg_ICACHE_TAG_WIDTH = 3;
									wire [2:0] icache_req_tag;
									// Trace: src/VX_fetch.sv:13:5
									wire icache_req_ready;
									// Trace: src/VX_fetch.sv:14:5
									wire [0:0] rsp_uuid;
									// Trace: src/VX_fetch.sv:15:5
									wire [1:0] req_tag;
									wire [1:0] rsp_tag;
									// Trace: src/VX_fetch.sv:16:5
									wire icache_req_fire = icache_req_valid && icache_req_ready;
									// Trace: src/VX_fetch.sv:17:5
									assign req_tag = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[35-:2];
									// Trace: src/VX_fetch.sv:18:5
									assign {rsp_uuid, rsp_tag} = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].rsp_data[2-:3];
									// Trace: src/VX_fetch.sv:19:5
									localparam VX_gpu_pkg_PC_BITS = 30;
									wire [29:0] rsp_PC;
									// Trace: src/VX_fetch.sv:20:5
									wire [3:0] rsp_tmask;
									// Trace: src/VX_fetch.sv:21:5
									VX_dp_ram #(
										.DATAW(34),
										.SIZE(4),
										.RDW_MODE("R"),
										.LUTRAM(1)
									) tag_store(
										.clk(clk),
										.reset(reset),
										.read(1'b1),
										.write(icache_req_fire),
										.wren(1'b1),
										.waddr(req_tag),
										.wdata({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[29-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[33-:4]}),
										.raddr(rsp_tag),
										.rdata({rsp_PC, rsp_tmask})
									);
									// Trace: src/VX_fetch.sv:37:5
									wire ibuf_ready = 1'b1;
									// Trace: src/VX_fetch.sv:38:5
									assign icache_req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.valid && ibuf_ready;
									// Trace: src/VX_fetch.sv:39:5
									assign icache_req_addr = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[0+:VX_gpu_pkg_ICACHE_ADDR_WIDTH];
									// Trace: src/VX_fetch.sv:40:5
									assign icache_req_tag = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.data[36-:1], req_tag};
									// Trace: src/VX_fetch.sv:41:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.schedule_if.ready = icache_req_ready && ibuf_ready;
									// Trace: src/VX_fetch.sv:42:5
									VX_elastic_buffer #(
										.DATAW(33),
										.SIZE(2),
										.OUT_REG(1)
									) req_buf(
										.clk(clk),
										.reset(reset),
										.valid_in(icache_req_valid),
										.ready_in(icache_req_ready),
										.data_in({icache_req_addr, icache_req_tag}),
										.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_data[71-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_data[2-:3]}),
										.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_valid),
										.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_ready)
									);
									// Trace: src/VX_fetch.sv:56:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_data[5-:3] = 1'sb0;
									// Trace: src/VX_fetch.sv:57:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_data[72] = 0;
									// Trace: src/VX_fetch.sv:58:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_data[9-:4] = 1'sb1;
									// Trace: src/VX_fetch.sv:59:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].req_data[41-:32] = 1'sb0;
									// Trace: src/VX_fetch.sv:60:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].rsp_valid;
									// Trace: src/VX_fetch.sv:61:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[65-:4] = rsp_tmask;
									// Trace: src/VX_fetch.sv:62:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[67-:2] = rsp_tag;
									// Trace: src/VX_fetch.sv:63:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[61-:30] = rsp_PC;
									// Trace: src/VX_fetch.sv:64:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[31-:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].rsp_data[34-:32];
									// Trace: src/VX_fetch.sv:65:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[68-:1] = rsp_uuid;
									// Trace: src/VX_fetch.sv:66:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_icache_bus_if[_mbase_icache_bus_if].rsp_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.ready;
								end
								assign fetch.clk = clk;
								assign fetch.reset = reset;
								// Trace: src/VX_core.sv:63:5
								// expanded module instance: decode
								localparam _param_21B54_INSTANCE_ID = "";
								if (1) begin : decode
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_decode.sv:2:15
									localparam INSTANCE_ID = _param_21B54_INSTANCE_ID;
									// Trace: src/VX_decode.sv:4:5
									wire clk;
									// Trace: src/VX_decode.sv:5:5
									wire reset;
									// Trace: src/VX_decode.sv:6:5
									// removed modport instance fetch_if
									// Trace: src/VX_decode.sv:7:5
									// removed modport instance decode_if
									// Trace: src/VX_decode.sv:8:5
									// removed modport instance decode_sched_if
									// Trace: src/VX_decode.sv:10:5
									localparam VX_gpu_pkg_EX_SFU = 2;
									localparam VX_gpu_pkg_EX_FPU = 2;
									localparam VX_gpu_pkg_EX_TCU = 2;
									localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
									localparam VX_gpu_pkg_EX_BITS = 2;
									localparam VX_gpu_pkg_INST_OP_BITS = 4;
									localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									localparam VX_gpu_pkg_PC_BITS = 30;
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
									// removed localparam type VX_gpu_pkg_alu_args_t
									localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
									// removed localparam type VX_gpu_pkg_csr_args_t
									localparam VX_gpu_pkg_INST_FMT_BITS = 2;
									localparam VX_gpu_pkg_INST_FRM_BITS = 3;
									// removed localparam type VX_gpu_pkg_fpu_args_t
									localparam VX_gpu_pkg_OFFSET_BITS = 12;
									// removed localparam type VX_gpu_pkg_lsu_args_t
									// removed localparam type VX_gpu_pkg_wctl_args_t
									// removed localparam type VX_gpu_pkg_op_args_t
									localparam VX_gpu_pkg_REG_TYPES = 1;
									localparam VX_gpu_pkg_REG_TYPE_BITS = 1;
									localparam VX_gpu_pkg_RV_REGS_BITS = 5;
									// removed localparam type VX_gpu_pkg_reg_idx_t
									// removed localparam type VX_gpu_pkg_decode_t
									localparam OUT_DATAW = 108;
									// Trace: src/VX_decode.sv:11:5
									reg [1:0] ex_type;
									// Trace: src/VX_decode.sv:12:5
									reg [3:0] op_type;
									// Trace: src/VX_decode.sv:13:5
									reg [36:0] op_args;
									// Trace: src/VX_decode.sv:14:5
									reg [5:0] rd_v;
									reg [5:0] rs1_v;
									reg [5:0] rs2_v;
									reg [5:0] rs3_v;
									// Trace: src/VX_decode.sv:15:5
									reg use_rd;
									reg use_rs1;
									reg use_rs2;
									reg use_rs3;
									// Trace: src/VX_decode.sv:16:5
									reg is_wstall;
									// Trace: src/VX_decode.sv:17:5
									wire [31:0] instr = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[31-:32];
									// Trace: src/VX_decode.sv:18:5
									wire [6:0] opcode = instr[6:0];
									// Trace: src/VX_decode.sv:19:5
									wire [1:0] funct2 = instr[26:25];
									// Trace: src/VX_decode.sv:20:5
									wire [2:0] funct3 = instr[14:12];
									// Trace: src/VX_decode.sv:21:5
									wire [4:0] funct5 = instr[31:27];
									// Trace: src/VX_decode.sv:22:5
									wire [6:0] funct7 = instr[31:25];
									// Trace: src/VX_decode.sv:23:5
									wire [11:0] u_12 = instr[31:20];
									// Trace: src/VX_decode.sv:24:5
									wire [4:0] rd = instr[11:7];
									// Trace: src/VX_decode.sv:25:5
									wire [4:0] rs1 = instr[19:15];
									// Trace: src/VX_decode.sv:26:5
									wire [4:0] rs2 = instr[24:20];
									// Trace: src/VX_decode.sv:27:5
									wire [4:0] rs3 = instr[31:27];
									// Trace: src/VX_decode.sv:28:5
									wire is_itype_sh = funct3[0] && ~funct3[1];
									// Trace: src/VX_decode.sv:29:5
									wire is_fpu_csr = u_12 <= 12'h003;
									// Trace: src/VX_decode.sv:30:5
									wire [19:0] ui_imm = instr[31:12];
									// Trace: src/VX_decode.sv:31:5
									wire [11:0] i_imm = (is_itype_sh ? {7'b0000000, instr[24:20]} : u_12);
									// Trace: src/VX_decode.sv:32:5
									wire [11:0] s_imm = {funct7, rd};
									// Trace: src/VX_decode.sv:33:5
									wire [12:0] b_imm = {instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};
									// Trace: src/VX_decode.sv:34:5
									wire [20:0] jal_imm = {instr[31], instr[19:12], instr[20], instr[30:21], 1'b0};
									// Trace: src/VX_decode.sv:35:5
									localparam VX_gpu_pkg_INST_ALU_BITS = 4;
									reg [3:0] r_type;
									// Trace: src/VX_decode.sv:36:5
									localparam VX_gpu_pkg_INST_ALU_ADD = 4'b0000;
									localparam VX_gpu_pkg_INST_ALU_AND = 4'b1100;
									localparam VX_gpu_pkg_INST_ALU_OR = 4'b1101;
									localparam VX_gpu_pkg_INST_ALU_SLL = 4'b1111;
									localparam VX_gpu_pkg_INST_ALU_SLT = 4'b0101;
									localparam VX_gpu_pkg_INST_ALU_SLTU = 4'b0100;
									localparam VX_gpu_pkg_INST_ALU_SRA = 4'b1001;
									localparam VX_gpu_pkg_INST_ALU_SRL = 4'b1000;
									localparam VX_gpu_pkg_INST_ALU_SUB = 4'b0111;
									localparam VX_gpu_pkg_INST_ALU_XOR = 4'b1110;
									always @(*)
										// Trace: src/VX_decode.sv:37:9
										case (funct3)
											3'h0:
												// Trace: src/VX_decode.sv:38:19
												r_type = (opcode[5] && funct7[5] ? VX_gpu_pkg_INST_ALU_SUB : VX_gpu_pkg_INST_ALU_ADD);
											3'h1:
												// Trace: src/VX_decode.sv:39:19
												r_type = VX_gpu_pkg_INST_ALU_SLL;
											3'h2:
												// Trace: src/VX_decode.sv:40:19
												r_type = VX_gpu_pkg_INST_ALU_SLT;
											3'h3:
												// Trace: src/VX_decode.sv:41:19
												r_type = VX_gpu_pkg_INST_ALU_SLTU;
											3'h4:
												// Trace: src/VX_decode.sv:42:19
												r_type = VX_gpu_pkg_INST_ALU_XOR;
											3'h5:
												// Trace: src/VX_decode.sv:43:19
												r_type = (funct7[5] ? VX_gpu_pkg_INST_ALU_SRA : VX_gpu_pkg_INST_ALU_SRL);
											3'h6:
												// Trace: src/VX_decode.sv:44:19
												r_type = VX_gpu_pkg_INST_ALU_OR;
											3'h7:
												// Trace: src/VX_decode.sv:45:19
												r_type = VX_gpu_pkg_INST_ALU_AND;
										endcase
									// Trace: src/VX_decode.sv:48:5
									localparam VX_gpu_pkg_INST_BR_BITS = 4;
									reg [3:0] b_type;
									// Trace: src/VX_decode.sv:49:5
									localparam VX_gpu_pkg_INST_BR_BEQ = 4'b0000;
									localparam VX_gpu_pkg_INST_BR_BGE = 4'b0111;
									localparam VX_gpu_pkg_INST_BR_BGEU = 4'b0110;
									localparam VX_gpu_pkg_INST_BR_BLT = 4'b0101;
									localparam VX_gpu_pkg_INST_BR_BLTU = 4'b0100;
									localparam VX_gpu_pkg_INST_BR_BNE = 4'b0010;
									always @(*)
										// Trace: src/VX_decode.sv:50:9
										case (funct3)
											3'h0:
												// Trace: src/VX_decode.sv:51:19
												b_type = VX_gpu_pkg_INST_BR_BEQ;
											3'h1:
												// Trace: src/VX_decode.sv:52:19
												b_type = VX_gpu_pkg_INST_BR_BNE;
											3'h4:
												// Trace: src/VX_decode.sv:53:19
												b_type = VX_gpu_pkg_INST_BR_BLT;
											3'h5:
												// Trace: src/VX_decode.sv:54:19
												b_type = VX_gpu_pkg_INST_BR_BGE;
											3'h6:
												// Trace: src/VX_decode.sv:55:19
												b_type = VX_gpu_pkg_INST_BR_BLTU;
											3'h7:
												// Trace: src/VX_decode.sv:56:19
												b_type = VX_gpu_pkg_INST_BR_BGEU;
											default:
												// Trace: src/VX_decode.sv:57:22
												b_type = 1'sbx;
										endcase
									// Trace: src/VX_decode.sv:60:5
									reg [3:0] s_type;
									// Trace: src/VX_decode.sv:61:5
									localparam VX_gpu_pkg_INST_BR_EBREAK = 4'b1011;
									localparam VX_gpu_pkg_INST_BR_ECALL = 4'b1010;
									localparam VX_gpu_pkg_INST_BR_MRET = 4'b1110;
									localparam VX_gpu_pkg_INST_BR_SRET = 4'b1101;
									localparam VX_gpu_pkg_INST_BR_URET = 4'b1100;
									always @(*)
										// Trace: src/VX_decode.sv:62:9
										case (u_12)
											12'h000:
												// Trace: src/VX_decode.sv:63:22
												s_type = VX_gpu_pkg_INST_BR_ECALL;
											12'h001:
												// Trace: src/VX_decode.sv:64:22
												s_type = VX_gpu_pkg_INST_BR_EBREAK;
											12'h002:
												// Trace: src/VX_decode.sv:65:22
												s_type = VX_gpu_pkg_INST_BR_URET;
											12'h102:
												// Trace: src/VX_decode.sv:66:22
												s_type = VX_gpu_pkg_INST_BR_SRET;
											12'h302:
												// Trace: src/VX_decode.sv:67:22
												s_type = VX_gpu_pkg_INST_BR_MRET;
											default:
												// Trace: src/VX_decode.sv:68:22
												s_type = 1'sbx;
										endcase
									// Trace: src/VX_decode.sv:71:5
									localparam VX_gpu_pkg_INST_M_BITS = 3;
									reg [2:0] m_type;
									// Trace: src/VX_decode.sv:72:5
									localparam VX_gpu_pkg_INST_M_DIV = 3'b100;
									localparam VX_gpu_pkg_INST_M_DIVU = 3'b101;
									localparam VX_gpu_pkg_INST_M_MUL = 3'b000;
									localparam VX_gpu_pkg_INST_M_MULH = 3'b010;
									localparam VX_gpu_pkg_INST_M_MULHSU = 3'b011;
									localparam VX_gpu_pkg_INST_M_MULHU = 3'b001;
									localparam VX_gpu_pkg_INST_M_REM = 3'b110;
									localparam VX_gpu_pkg_INST_M_REMU = 3'b111;
									always @(*)
										// Trace: src/VX_decode.sv:73:9
										case (funct3)
											3'h0:
												// Trace: src/VX_decode.sv:74:19
												m_type = VX_gpu_pkg_INST_M_MUL;
											3'h1:
												// Trace: src/VX_decode.sv:75:19
												m_type = VX_gpu_pkg_INST_M_MULH;
											3'h2:
												// Trace: src/VX_decode.sv:76:19
												m_type = VX_gpu_pkg_INST_M_MULHSU;
											3'h3:
												// Trace: src/VX_decode.sv:77:19
												m_type = VX_gpu_pkg_INST_M_MULHU;
											3'h4:
												// Trace: src/VX_decode.sv:78:19
												m_type = VX_gpu_pkg_INST_M_DIV;
											3'h5:
												// Trace: src/VX_decode.sv:79:19
												m_type = VX_gpu_pkg_INST_M_DIVU;
											3'h6:
												// Trace: src/VX_decode.sv:80:19
												m_type = VX_gpu_pkg_INST_M_REM;
											3'h7:
												// Trace: src/VX_decode.sv:81:19
												m_type = VX_gpu_pkg_INST_M_REMU;
										endcase
									// Trace: src/VX_decode.sv:84:5
									localparam VX_gpu_pkg_ALU_TYPE_ARITH = 0;
									localparam VX_gpu_pkg_ALU_TYPE_BRANCH = 1;
									localparam VX_gpu_pkg_ALU_TYPE_MULDIV = 2;
									localparam VX_gpu_pkg_ALU_TYPE_OTHER = 3;
									localparam VX_gpu_pkg_EX_ALU = 0;
									localparam VX_gpu_pkg_EX_LSU = 1;
									localparam VX_gpu_pkg_INST_ALU_AUIPC = 4'b0011;
									localparam VX_gpu_pkg_INST_ALU_CZEQ = 4'b1010;
									localparam VX_gpu_pkg_INST_ALU_CZNE = 4'b1011;
									localparam VX_gpu_pkg_INST_ALU_LUI = 4'b0010;
									localparam VX_gpu_pkg_INST_AUIPC = 7'b0010111;
									localparam VX_gpu_pkg_INST_B = 7'b1100011;
									localparam VX_gpu_pkg_INST_BR_JAL = 4'b1000;
									localparam VX_gpu_pkg_INST_BR_JALR = 4'b1001;
									localparam VX_gpu_pkg_INST_EXT1 = 7'b0001011;
									localparam VX_gpu_pkg_INST_FENCE = 7'b0001111;
									localparam VX_gpu_pkg_INST_I = 7'b0010011;
									localparam VX_gpu_pkg_INST_JAL = 7'b1101111;
									localparam VX_gpu_pkg_INST_JALR = 7'b1100111;
									localparam VX_gpu_pkg_INST_L = 7'b0000011;
									localparam VX_gpu_pkg_INST_LSU_FENCE = 4'b1111;
									localparam VX_gpu_pkg_INST_LUI = 7'b0110111;
									localparam VX_gpu_pkg_INST_R = 7'b0110011;
									localparam VX_gpu_pkg_INST_R_F7_MUL = 7'b0000001;
									localparam VX_gpu_pkg_INST_R_F7_ZICOND = 7'b0000111;
									localparam VX_gpu_pkg_INST_S = 7'b0100011;
									localparam VX_gpu_pkg_INST_SFU_BAR = 4'h4;
									localparam VX_gpu_pkg_INST_SFU_JOIN = 4'h3;
									localparam VX_gpu_pkg_INST_SFU_PRED = 4'h5;
									localparam VX_gpu_pkg_INST_SFU_SPLIT = 4'h2;
									localparam VX_gpu_pkg_INST_SFU_TMC = 4'h0;
									localparam VX_gpu_pkg_INST_SFU_WSPAWN = 4'h1;
									localparam VX_gpu_pkg_INST_SYS = 7'b1110011;
									function automatic [3:0] VX_gpu_pkg_inst_sfu_csr;
										// Trace: src/VX_gpu_pkg.sv:249:49
										input reg [2:0] funct3;
										// Trace: src/VX_gpu_pkg.sv:250:9
										VX_gpu_pkg_inst_sfu_csr = (4'h6 + sv2v_cast_4(funct3[1:0])) - 4'h1;
									endfunction
									always @(*) begin
										// Trace: src/VX_decode.sv:85:9
										ex_type = 1'sbx;
										// Trace: src/VX_decode.sv:86:9
										op_type = 1'sbx;
										// Trace: src/VX_decode.sv:87:9
										op_args = 1'sbx;
										// Trace: src/VX_decode.sv:88:9
										rd_v = 1'sbx;
										// Trace: src/VX_decode.sv:89:9
										rs1_v = 1'sbx;
										// Trace: src/VX_decode.sv:90:9
										rs2_v = 1'sbx;
										// Trace: src/VX_decode.sv:91:9
										rs3_v = 1'sbx;
										// Trace: src/VX_decode.sv:92:9
										use_rd = 0;
										// Trace: src/VX_decode.sv:93:9
										use_rs1 = 0;
										// Trace: src/VX_decode.sv:94:9
										use_rs2 = 0;
										// Trace: src/VX_decode.sv:95:9
										use_rs3 = 0;
										// Trace: src/VX_decode.sv:96:9
										is_wstall = 0;
										// Trace: src/VX_decode.sv:97:9
										case (opcode)
											VX_gpu_pkg_INST_I: begin
												// Trace: src/VX_decode.sv:99:17
												ex_type = VX_gpu_pkg_EX_ALU;
												// Trace: src/VX_decode.sv:100:17
												op_type = r_type;
												// Trace: src/VX_decode.sv:101:17
												op_args[33-:2] = VX_gpu_pkg_ALU_TYPE_ARITH;
												// Trace: src/VX_decode.sv:102:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:103:17
												op_args[36] = 0;
												// Trace: src/VX_decode.sv:104:17
												op_args[35] = 1;
												// Trace: src/VX_decode.sv:105:17
												op_args[31-:32] = {{21 {i_imm[11]}}, i_imm[10:0]};
												// Trace: src/VX_decode.sv:106:5
												rd_v[4-:5] = rd;
												// Trace: src/VX_decode.sv:107:5
												rd_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:108:5
												use_rd = 1;
												// Trace: src/VX_decode.sv:109:5
												rs1_v[4-:5] = rs1;
												// Trace: src/VX_decode.sv:110:5
												rs1_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:111:5
												use_rs1 = 1;
											end
											VX_gpu_pkg_INST_R: begin
												// Trace: src/VX_decode.sv:114:17
												ex_type = VX_gpu_pkg_EX_ALU;
												// Trace: src/VX_decode.sv:115:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:116:17
												op_args[36] = 0;
												// Trace: src/VX_decode.sv:117:17
												op_args[35] = 0;
												// Trace: src/VX_decode.sv:118:5
												rd_v[4-:5] = rd;
												// Trace: src/VX_decode.sv:119:5
												rd_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:120:5
												use_rd = 1;
												// Trace: src/VX_decode.sv:121:5
												rs1_v[4-:5] = rs1;
												// Trace: src/VX_decode.sv:122:5
												rs1_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:123:5
												use_rs1 = 1;
												// Trace: src/VX_decode.sv:124:5
												rs2_v[4-:5] = rs2;
												// Trace: src/VX_decode.sv:125:5
												rs2_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:126:5
												use_rs2 = 1;
												// Trace: src/VX_decode.sv:127:17
												case (funct7)
													VX_gpu_pkg_INST_R_F7_MUL: begin
														// Trace: src/VX_decode.sv:129:25
														op_type = sv2v_cast_4(m_type);
														// Trace: src/VX_decode.sv:130:25
														op_args[33-:2] = VX_gpu_pkg_ALU_TYPE_MULDIV;
													end
													VX_gpu_pkg_INST_R_F7_ZICOND: begin
														// Trace: src/VX_decode.sv:133:25
														op_type = (funct3[1] ? VX_gpu_pkg_INST_ALU_CZNE : VX_gpu_pkg_INST_ALU_CZEQ);
														// Trace: src/VX_decode.sv:134:25
														op_args[33-:2] = VX_gpu_pkg_ALU_TYPE_ARITH;
													end
													default: begin
														// Trace: src/VX_decode.sv:137:25
														op_type = r_type;
														// Trace: src/VX_decode.sv:138:25
														op_args[33-:2] = VX_gpu_pkg_ALU_TYPE_ARITH;
													end
												endcase
											end
											VX_gpu_pkg_INST_LUI: begin
												// Trace: src/VX_decode.sv:143:17
												ex_type = VX_gpu_pkg_EX_ALU;
												// Trace: src/VX_decode.sv:144:17
												op_type = VX_gpu_pkg_INST_ALU_LUI;
												// Trace: src/VX_decode.sv:145:17
												op_args[33-:2] = VX_gpu_pkg_ALU_TYPE_ARITH;
												// Trace: src/VX_decode.sv:146:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:147:17
												op_args[36] = 0;
												// Trace: src/VX_decode.sv:148:17
												op_args[35] = 1;
												// Trace: src/VX_decode.sv:149:17
												op_args[31-:32] = {ui_imm[19], ui_imm[18:0], 12'sd0};
												// Trace: src/VX_decode.sv:150:5
												rd_v[4-:5] = rd;
												// Trace: src/VX_decode.sv:151:5
												rd_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:152:5
												use_rd = 1;
											end
											VX_gpu_pkg_INST_AUIPC: begin
												// Trace: src/VX_decode.sv:155:17
												ex_type = VX_gpu_pkg_EX_ALU;
												// Trace: src/VX_decode.sv:156:17
												op_type = VX_gpu_pkg_INST_ALU_AUIPC;
												// Trace: src/VX_decode.sv:157:17
												op_args[33-:2] = VX_gpu_pkg_ALU_TYPE_ARITH;
												// Trace: src/VX_decode.sv:158:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:159:17
												op_args[36] = 1;
												// Trace: src/VX_decode.sv:160:17
												op_args[35] = 1;
												// Trace: src/VX_decode.sv:161:17
												op_args[31-:32] = {ui_imm[19], ui_imm[18:0], 12'sd0};
												// Trace: src/VX_decode.sv:162:5
												rd_v[4-:5] = rd;
												// Trace: src/VX_decode.sv:163:5
												rd_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:164:5
												use_rd = 1;
											end
											VX_gpu_pkg_INST_JAL: begin
												// Trace: src/VX_decode.sv:167:17
												ex_type = VX_gpu_pkg_EX_ALU;
												// Trace: src/VX_decode.sv:168:17
												op_type = VX_gpu_pkg_INST_BR_JAL;
												// Trace: src/VX_decode.sv:169:17
												op_args[33-:2] = VX_gpu_pkg_ALU_TYPE_BRANCH;
												// Trace: src/VX_decode.sv:170:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:171:17
												op_args[36] = 1;
												// Trace: src/VX_decode.sv:172:17
												op_args[35] = 1;
												// Trace: src/VX_decode.sv:173:17
												op_args[31-:32] = {{12 {jal_imm[20]}}, jal_imm[19:0]};
												// Trace: src/VX_decode.sv:174:17
												is_wstall = 1;
												// Trace: src/VX_decode.sv:175:5
												rd_v[4-:5] = rd;
												// Trace: src/VX_decode.sv:176:5
												rd_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:177:5
												use_rd = 1;
											end
											VX_gpu_pkg_INST_JALR: begin
												// Trace: src/VX_decode.sv:180:17
												ex_type = VX_gpu_pkg_EX_ALU;
												// Trace: src/VX_decode.sv:181:17
												op_type = VX_gpu_pkg_INST_BR_JALR;
												// Trace: src/VX_decode.sv:182:17
												op_args[33-:2] = VX_gpu_pkg_ALU_TYPE_BRANCH;
												// Trace: src/VX_decode.sv:183:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:184:17
												op_args[36] = 0;
												// Trace: src/VX_decode.sv:185:17
												op_args[35] = 1;
												// Trace: src/VX_decode.sv:186:17
												op_args[31-:32] = {{21 {u_12[11]}}, u_12[10:0]};
												// Trace: src/VX_decode.sv:187:17
												is_wstall = 1;
												// Trace: src/VX_decode.sv:188:5
												rd_v[4-:5] = rd;
												// Trace: src/VX_decode.sv:189:5
												rd_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:190:5
												use_rd = 1;
												// Trace: src/VX_decode.sv:191:5
												rs1_v[4-:5] = rs1;
												// Trace: src/VX_decode.sv:192:5
												rs1_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:193:5
												use_rs1 = 1;
											end
											VX_gpu_pkg_INST_B: begin
												// Trace: src/VX_decode.sv:196:17
												ex_type = VX_gpu_pkg_EX_ALU;
												// Trace: src/VX_decode.sv:197:17
												op_type = b_type;
												// Trace: src/VX_decode.sv:198:17
												op_args[33-:2] = VX_gpu_pkg_ALU_TYPE_BRANCH;
												// Trace: src/VX_decode.sv:199:17
												op_args[34] = 0;
												// Trace: src/VX_decode.sv:200:17
												op_args[36] = 1;
												// Trace: src/VX_decode.sv:201:17
												op_args[35] = 1;
												// Trace: src/VX_decode.sv:202:17
												op_args[31-:32] = {{20 {b_imm[12]}}, b_imm[11:0]};
												// Trace: src/VX_decode.sv:203:17
												is_wstall = 1;
												// Trace: src/VX_decode.sv:204:5
												rs1_v[4-:5] = rs1;
												// Trace: src/VX_decode.sv:205:5
												rs1_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:206:5
												use_rs1 = 1;
												// Trace: src/VX_decode.sv:207:5
												rs2_v[4-:5] = rs2;
												// Trace: src/VX_decode.sv:208:5
												rs2_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:209:5
												use_rs2 = 1;
											end
											VX_gpu_pkg_INST_FENCE: begin
												// Trace: src/VX_decode.sv:212:17
												ex_type = VX_gpu_pkg_EX_LSU;
												// Trace: src/VX_decode.sv:213:17
												op_type = VX_gpu_pkg_INST_LSU_FENCE;
												// Trace: src/VX_decode.sv:214:17
												op_args[13] = 0;
												// Trace: src/VX_decode.sv:215:17
												op_args[12] = 0;
												// Trace: src/VX_decode.sv:216:17
												op_args[11-:12] = 0;
											end
											VX_gpu_pkg_INST_SYS:
												// Trace: src/VX_decode.sv:219:17
												if (funct3[1:0] != 0) begin
													// Trace: src/VX_decode.sv:220:21
													ex_type = VX_gpu_pkg_EX_SFU;
													// Trace: src/VX_decode.sv:221:21
													op_type = VX_gpu_pkg_inst_sfu_csr(funct3);
													// Trace: src/VX_decode.sv:222:21
													op_args[16-:12] = u_12;
													// Trace: src/VX_decode.sv:223:21
													op_args[17] = funct3[2];
													// Trace: src/VX_decode.sv:224:21
													is_wstall = is_fpu_csr;
													// Trace: src/VX_decode.sv:225:5
													rd_v[4-:5] = rd;
													// Trace: src/VX_decode.sv:226:5
													rd_v[5-:1] = 0;
													// Trace: src/VX_decode.sv:227:5
													use_rd = 1;
													// Trace: src/VX_decode.sv:228:21
													if (funct3[2])
														// Trace: src/VX_decode.sv:229:25
														op_args[4-:5] = rs1;
													else begin
														// Trace: src/VX_decode.sv:231:5
														rs1_v[4-:5] = rs1;
														// Trace: src/VX_decode.sv:232:5
														rs1_v[5-:1] = 0;
														// Trace: src/VX_decode.sv:233:5
														use_rs1 = 1;
													end
												end
												else begin
													// Trace: src/VX_decode.sv:236:21
													ex_type = VX_gpu_pkg_EX_ALU;
													// Trace: src/VX_decode.sv:237:21
													op_type = s_type;
													// Trace: src/VX_decode.sv:238:21
													op_args[33-:2] = VX_gpu_pkg_ALU_TYPE_BRANCH;
													// Trace: src/VX_decode.sv:239:21
													op_args[34] = 0;
													// Trace: src/VX_decode.sv:240:21
													op_args[35] = 1;
													// Trace: src/VX_decode.sv:241:21
													op_args[36] = 1;
													// Trace: src/VX_decode.sv:242:21
													op_args[31-:32] = 32'd4;
													// Trace: src/VX_decode.sv:243:21
													is_wstall = 1;
													// Trace: src/VX_decode.sv:244:5
													rd_v[4-:5] = rd;
													// Trace: src/VX_decode.sv:245:5
													rd_v[5-:1] = 0;
													// Trace: src/VX_decode.sv:246:5
													use_rd = 1;
												end
											VX_gpu_pkg_INST_L: begin
												// Trace: src/VX_decode.sv:250:17
												ex_type = VX_gpu_pkg_EX_LSU;
												// Trace: src/VX_decode.sv:251:17
												op_type = sv2v_cast_4({1'b0, funct3});
												// Trace: src/VX_decode.sv:252:17
												op_args[13] = 0;
												// Trace: src/VX_decode.sv:253:17
												op_args[12] = opcode[2];
												// Trace: src/VX_decode.sv:254:17
												op_args[11-:12] = u_12;
												// Trace: src/VX_decode.sv:255:5
												rs1_v[4-:5] = rs1;
												// Trace: src/VX_decode.sv:256:5
												rs1_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:257:5
												use_rs1 = 1;
												// Trace: src/VX_decode.sv:258:5
												rd_v[4-:5] = rd;
												// Trace: src/VX_decode.sv:259:5
												rd_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:260:5
												use_rd = 1;
											end
											VX_gpu_pkg_INST_S: begin
												// Trace: src/VX_decode.sv:263:17
												ex_type = VX_gpu_pkg_EX_LSU;
												// Trace: src/VX_decode.sv:264:17
												op_type = sv2v_cast_4({1'b1, funct3});
												// Trace: src/VX_decode.sv:265:17
												op_args[13] = 1;
												// Trace: src/VX_decode.sv:266:17
												op_args[12] = opcode[2];
												// Trace: src/VX_decode.sv:267:17
												op_args[11-:12] = s_imm;
												// Trace: src/VX_decode.sv:268:5
												rs1_v[4-:5] = rs1;
												// Trace: src/VX_decode.sv:269:5
												rs1_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:270:5
												use_rs1 = 1;
												// Trace: src/VX_decode.sv:271:5
												rs2_v[4-:5] = rs2;
												// Trace: src/VX_decode.sv:272:5
												rs2_v[5-:1] = 0;
												// Trace: src/VX_decode.sv:273:5
												use_rs2 = 1;
											end
											VX_gpu_pkg_INST_EXT1:
												// Trace: src/VX_decode.sv:276:17
												case (funct7)
													7'h00: begin
														// Trace: src/VX_decode.sv:278:25
														ex_type = VX_gpu_pkg_EX_SFU;
														// Trace: src/VX_decode.sv:279:25
														is_wstall = 1;
														// Trace: src/VX_decode.sv:280:25
														case (funct3)
															3'h0: begin
																// Trace: src/VX_decode.sv:282:33
																op_type = VX_gpu_pkg_INST_SFU_TMC;
																// Trace: src/VX_decode.sv:283:5
																rs1_v[4-:5] = rs1;
																// Trace: src/VX_decode.sv:284:5
																rs1_v[5-:1] = 0;
																// Trace: src/VX_decode.sv:285:5
																use_rs1 = 1;
															end
															3'h1: begin
																// Trace: src/VX_decode.sv:288:33
																op_type = VX_gpu_pkg_INST_SFU_WSPAWN;
																// Trace: src/VX_decode.sv:289:5
																rs1_v[4-:5] = rs1;
																// Trace: src/VX_decode.sv:290:5
																rs1_v[5-:1] = 0;
																// Trace: src/VX_decode.sv:291:5
																use_rs1 = 1;
																// Trace: src/VX_decode.sv:292:5
																rs2_v[4-:5] = rs2;
																// Trace: src/VX_decode.sv:293:5
																rs2_v[5-:1] = 0;
																// Trace: src/VX_decode.sv:294:5
																use_rs2 = 1;
															end
															3'h2: begin
																// Trace: src/VX_decode.sv:297:33
																op_type = VX_gpu_pkg_INST_SFU_SPLIT;
																// Trace: src/VX_decode.sv:298:33
																op_args[0] = rs2[0];
																// Trace: src/VX_decode.sv:299:5
																rs1_v[4-:5] = rs1;
																// Trace: src/VX_decode.sv:300:5
																rs1_v[5-:1] = 0;
																// Trace: src/VX_decode.sv:301:5
																use_rs1 = 1;
																// Trace: src/VX_decode.sv:302:5
																rd_v[4-:5] = rd;
																// Trace: src/VX_decode.sv:303:5
																rd_v[5-:1] = 0;
																// Trace: src/VX_decode.sv:304:5
																use_rd = 1;
															end
															3'h3: begin
																// Trace: src/VX_decode.sv:307:33
																op_type = VX_gpu_pkg_INST_SFU_JOIN;
																// Trace: src/VX_decode.sv:308:5
																rs1_v[4-:5] = rs1;
																// Trace: src/VX_decode.sv:309:5
																rs1_v[5-:1] = 0;
																// Trace: src/VX_decode.sv:310:5
																use_rs1 = 1;
															end
															3'h4: begin
																// Trace: src/VX_decode.sv:313:33
																op_type = VX_gpu_pkg_INST_SFU_BAR;
																// Trace: src/VX_decode.sv:314:5
																rs1_v[4-:5] = rs1;
																// Trace: src/VX_decode.sv:315:5
																rs1_v[5-:1] = 0;
																// Trace: src/VX_decode.sv:316:5
																use_rs1 = 1;
																// Trace: src/VX_decode.sv:317:5
																rs2_v[4-:5] = rs2;
																// Trace: src/VX_decode.sv:318:5
																rs2_v[5-:1] = 0;
																// Trace: src/VX_decode.sv:319:5
																use_rs2 = 1;
															end
															3'h5: begin
																// Trace: src/VX_decode.sv:322:33
																op_type = VX_gpu_pkg_INST_SFU_PRED;
																// Trace: src/VX_decode.sv:323:33
																op_args[0] = rd[0];
																// Trace: src/VX_decode.sv:324:5
																rs1_v[4-:5] = rs1;
																// Trace: src/VX_decode.sv:325:5
																rs1_v[5-:1] = 0;
																// Trace: src/VX_decode.sv:326:5
																use_rs1 = 1;
																// Trace: src/VX_decode.sv:327:5
																rs2_v[4-:5] = rs2;
																// Trace: src/VX_decode.sv:328:5
																rs2_v[5-:1] = 0;
																// Trace: src/VX_decode.sv:329:5
																use_rs2 = 1;
															end
															default:
																;
														endcase
													end
													7'h01: begin
														// Trace: src/VX_decode.sv:335:25
														ex_type = VX_gpu_pkg_EX_ALU;
														// Trace: src/VX_decode.sv:336:25
														op_args[33-:2] = VX_gpu_pkg_ALU_TYPE_OTHER;
														// Trace: src/VX_decode.sv:337:25
														use_rd = 1;
														// Trace: src/VX_decode.sv:338:5
														rd_v[4-:5] = rd;
														// Trace: src/VX_decode.sv:339:5
														rd_v[5-:1] = 0;
														// Trace: src/VX_decode.sv:340:5
														use_rd = 1;
														// Trace: src/VX_decode.sv:341:5
														rs1_v[4-:5] = rs1;
														// Trace: src/VX_decode.sv:342:5
														rs1_v[5-:1] = 0;
														// Trace: src/VX_decode.sv:343:5
														use_rs1 = 1;
														// Trace: src/VX_decode.sv:344:25
														if (funct3[2]) begin
															// Trace: src/VX_decode.sv:345:5
															rs2_v[4-:5] = rs2;
															// Trace: src/VX_decode.sv:346:5
															rs2_v[5-:1] = 0;
															// Trace: src/VX_decode.sv:347:5
															use_rs2 = 1;
														end
														// Trace: src/VX_decode.sv:349:25
														op_type = sv2v_cast_4(funct3);
													end
													default:
														;
												endcase
											default:
												;
										endcase
									end
									// Trace: src/VX_decode.sv:357:5
									wire wb = use_rd && (rd_v != 0);
									// Trace: src/VX_decode.sv:358:5
									wire [2:0] used_rs = {use_rs3, use_rs2, use_rs1};
									// Trace: src/VX_decode.sv:359:5
									VX_elastic_buffer #(
										.DATAW(OUT_DATAW),
										.SIZE(0)
									) req_buf(
										.clk(clk),
										.reset(reset),
										.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.valid),
										.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.ready),
										.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[68-:1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[67-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[65-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[61-:30], ex_type, op_type, op_args, wb, used_rs, rd_v, rs1_v, rs2_v, rs3_v}),
										.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[107], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[106-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[104-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[100-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[70-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[68-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[64-:37], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[27], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[26-:3], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[23-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[17-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[11-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[5-:6]}),
										.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.valid),
										.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.ready)
									);
									// Trace: src/VX_decode.sv:372:5
									wire fetch_fire = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.ready;
									// Trace: src/VX_decode.sv:373:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.valid = fetch_fire;
									// Trace: src/VX_decode.sv:374:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.fetch_if.data[67-:2];
									// Trace: src/VX_decode.sv:375:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_sched_if.unlock = ~is_wstall;
								end
								assign decode.clk = clk;
								assign decode.reset = reset;
								// Trace: src/VX_core.sv:72:5
								// expanded module instance: issue
								localparam _bbase_CF65A_writeback_if = 0;
								localparam _bbase_CF65A_dispatch_if = 0;
								localparam _bbase_CF65A_issue_sched_if = 0;
								localparam _param_CF65A_INSTANCE_ID = "";
								if (1) begin : issue
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_issue.sv:2:15
									localparam INSTANCE_ID = _param_CF65A_INSTANCE_ID;
									// Trace: src/VX_issue.sv:4:5
									wire clk;
									// Trace: src/VX_issue.sv:5:5
									wire reset;
									// Trace: src/VX_issue.sv:6:5
									// removed modport instance decode_if
									// Trace: src/VX_issue.sv:7:5
									localparam _mbase_writeback_if = 0;
									// Trace: src/VX_issue.sv:8:5
									localparam VX_gpu_pkg_EX_SFU = 2;
									localparam VX_gpu_pkg_EX_FPU = 2;
									localparam VX_gpu_pkg_EX_TCU = 2;
									localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
									localparam _mbase_dispatch_if = 0;
									// Trace: src/VX_issue.sv:9:5
									localparam _mbase_issue_sched_if = 0;
									// Trace: src/VX_issue.sv:11:5
									localparam VX_gpu_pkg_ISSUE_ISW_BITS = 0;
									localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									function automatic [0:0] VX_gpu_pkg_wid_to_isw;
										// Trace: src/VX_gpu_pkg.sv:276:9
										input reg [1:0] wid;
										// Trace: src/VX_gpu_pkg.sv:278:9
										begin
											// Trace: src/VX_gpu_pkg.sv:281:13
											VX_gpu_pkg_wid_to_isw = 0;
										end
									endfunction
									wire [0:0] decode_isw = VX_gpu_pkg_wid_to_isw(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data[106-:2]);
									// Trace: src/VX_issue.sv:12:5
									wire [0:0] decode_ready_in;
									// Trace: src/VX_issue.sv:13:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.ready = decode_ready_in[decode_isw];
									// Trace: src/VX_issue.sv:15:5
									genvar _gv_issue_id_1;
									for (_gv_issue_id_1 = 0; _gv_issue_id_1 < 1; _gv_issue_id_1 = _gv_issue_id_1 + 1) begin : g_slices
										localparam issue_id = _gv_issue_id_1;
										// Trace: src/VX_issue.sv:16:9
										// expanded interface instance: slice_decode_if
										if (1) begin : slice_decode_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_decode_if.sv:2:5
											wire valid;
											// Trace: src/VX_decode_if.sv:3:5
											localparam VX_gpu_pkg_EX_SFU = 2;
											localparam VX_gpu_pkg_EX_FPU = 2;
											localparam VX_gpu_pkg_EX_TCU = 2;
											localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
											localparam VX_gpu_pkg_EX_BITS = 2;
											localparam VX_gpu_pkg_INST_OP_BITS = 4;
											localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
											// removed localparam type VX_gpu_pkg_alu_args_t
											localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
											// removed localparam type VX_gpu_pkg_csr_args_t
											localparam VX_gpu_pkg_INST_FMT_BITS = 2;
											localparam VX_gpu_pkg_INST_FRM_BITS = 3;
											// removed localparam type VX_gpu_pkg_fpu_args_t
											localparam VX_gpu_pkg_OFFSET_BITS = 12;
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_REG_TYPE_BITS = 1;
											localparam VX_gpu_pkg_RV_REGS_BITS = 5;
											// removed localparam type VX_gpu_pkg_reg_idx_t
											// removed localparam type VX_gpu_pkg_decode_t
											wire [107:0] data;
											// Trace: src/VX_decode_if.sv:4:5
											wire ready;
											// Trace: src/VX_decode_if.sv:5:5
											// Trace: src/VX_decode_if.sv:10:5
										end
										// Trace: src/VX_issue.sv:17:9
										// expanded interface instance: per_issue_dispatch_if
										genvar _arr_18544;
										for (_arr_18544 = 0; _arr_18544 <= 2; _arr_18544 = _arr_18544 + 1) begin : per_issue_dispatch_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_dispatch_if.sv:2:5
											wire valid;
											// Trace: src/VX_dispatch_if.sv:3:5
											localparam VX_gpu_pkg_INST_ALU_BITS = 4;
											localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
											localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
											localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_SIMD_COUNT = 1;
											localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
											localparam VX_gpu_pkg_SIMD_IDX_W = 1;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
											// removed localparam type VX_gpu_pkg_alu_args_t
											localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
											// removed localparam type VX_gpu_pkg_csr_args_t
											localparam VX_gpu_pkg_INST_FMT_BITS = 2;
											localparam VX_gpu_pkg_INST_FRM_BITS = 3;
											// removed localparam type VX_gpu_pkg_fpu_args_t
											localparam VX_gpu_pkg_OFFSET_BITS = 12;
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											// removed localparam type VX_gpu_pkg_dispatch_t
											wire [470:0] data;
											// Trace: src/VX_dispatch_if.sv:4:5
											wire ready;
											// Trace: src/VX_dispatch_if.sv:5:5
											// Trace: src/VX_dispatch_if.sv:10:5
										end
										// Trace: src/VX_issue.sv:18:9
										assign slice_decode_if.valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.valid && (decode_isw == issue_id);
										// Trace: src/VX_issue.sv:19:9
										assign slice_decode_if.data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.decode_if.data;
										// Trace: src/VX_issue.sv:20:9
										assign decode_ready_in[issue_id] = slice_decode_if.ready;
										// Trace: src/VX_issue.sv:21:9
										// expanded module instance: issue_slice
										localparam _bbase_A8822_writeback_if = issue_id + _mbase_writeback_if;
										localparam _bbase_A8822_dispatch_if = 0;
										localparam _bbase_A8822_issue_sched_if = issue_id + _mbase_issue_sched_if;
										localparam _param_A8822_INSTANCE_ID = "";
										localparam _param_A8822_ISSUE_ID = issue_id;
										if (1) begin : issue_slice
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_issue_slice.sv:2:15
											localparam INSTANCE_ID = _param_A8822_INSTANCE_ID;
											// Trace: src/VX_issue_slice.sv:3:15
											localparam ISSUE_ID = _param_A8822_ISSUE_ID;
											// Trace: src/VX_issue_slice.sv:5:5
											wire clk;
											// Trace: src/VX_issue_slice.sv:6:5
											wire reset;
											// Trace: src/VX_issue_slice.sv:7:5
											// removed modport instance decode_if
											// Trace: src/VX_issue_slice.sv:8:5
											localparam _mbase_writeback_if = _bbase_A8822_writeback_if;
											// Trace: src/VX_issue_slice.sv:9:5
											localparam VX_gpu_pkg_EX_SFU = 2;
											localparam VX_gpu_pkg_EX_FPU = 2;
											localparam VX_gpu_pkg_EX_TCU = 2;
											localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
											localparam _mbase_dispatch_if = 0;
											// Trace: src/VX_issue_slice.sv:10:5
											localparam _mbase_issue_sched_if = _bbase_A8822_issue_sched_if;
											// Trace: src/VX_issue_slice.sv:12:5
											localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
											// expanded interface instance: ibuffer_if
											genvar _arr_F0EBA;
											for (_arr_F0EBA = 0; _arr_F0EBA <= 3; _arr_F0EBA = _arr_F0EBA + 1) begin : ibuffer_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_ibuffer_if.sv:2:5
												wire valid;
												// Trace: src/VX_ibuffer_if.sv:3:5
												localparam VX_gpu_pkg_EX_SFU = 2;
												localparam VX_gpu_pkg_EX_FPU = 2;
												localparam VX_gpu_pkg_EX_TCU = 2;
												localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
												localparam VX_gpu_pkg_EX_BITS = 2;
												localparam VX_gpu_pkg_INST_OP_BITS = 4;
												localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
												localparam VX_gpu_pkg_PC_BITS = 30;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
												// removed localparam type VX_gpu_pkg_alu_args_t
												localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
												// removed localparam type VX_gpu_pkg_csr_args_t
												localparam VX_gpu_pkg_INST_FMT_BITS = 2;
												localparam VX_gpu_pkg_INST_FRM_BITS = 3;
												// removed localparam type VX_gpu_pkg_fpu_args_t
												localparam VX_gpu_pkg_OFFSET_BITS = 12;
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_REG_TYPE_BITS = 1;
												localparam VX_gpu_pkg_RV_REGS_BITS = 5;
												// removed localparam type VX_gpu_pkg_reg_idx_t
												// removed localparam type VX_gpu_pkg_ibuffer_t
												wire [105:0] data;
												// Trace: src/VX_ibuffer_if.sv:4:5
												wire ready;
												// Trace: src/VX_ibuffer_if.sv:5:5
												// Trace: src/VX_ibuffer_if.sv:10:5
											end
											// Trace: src/VX_issue_slice.sv:13:5
											// expanded interface instance: scoreboard_if
											if (1) begin : scoreboard_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_scoreboard_if.sv:2:5
												wire valid;
												// Trace: src/VX_scoreboard_if.sv:3:5
												localparam VX_gpu_pkg_EX_SFU = 2;
												localparam VX_gpu_pkg_EX_FPU = 2;
												localparam VX_gpu_pkg_EX_TCU = 2;
												localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
												localparam VX_gpu_pkg_EX_BITS = 2;
												localparam VX_gpu_pkg_INST_OP_BITS = 4;
												localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
												localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
												localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
												localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
												localparam VX_gpu_pkg_PC_BITS = 30;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
												// removed localparam type VX_gpu_pkg_alu_args_t
												localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
												// removed localparam type VX_gpu_pkg_csr_args_t
												localparam VX_gpu_pkg_INST_FMT_BITS = 2;
												localparam VX_gpu_pkg_INST_FRM_BITS = 3;
												// removed localparam type VX_gpu_pkg_fpu_args_t
												localparam VX_gpu_pkg_OFFSET_BITS = 12;
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_REG_TYPE_BITS = 1;
												localparam VX_gpu_pkg_RV_REGS_BITS = 5;
												// removed localparam type VX_gpu_pkg_reg_idx_t
												// removed localparam type VX_gpu_pkg_scoreboard_t
												wire [107:0] data;
												// Trace: src/VX_scoreboard_if.sv:4:5
												wire ready;
												// Trace: src/VX_scoreboard_if.sv:5:5
												// Trace: src/VX_scoreboard_if.sv:10:5
											end
											// Trace: src/VX_issue_slice.sv:14:5
											// expanded interface instance: operands_if
											if (1) begin : operands_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_operands_if.sv:2:5
												wire valid;
												// Trace: src/VX_operands_if.sv:3:5
												localparam VX_gpu_pkg_EX_SFU = 2;
												localparam VX_gpu_pkg_EX_FPU = 2;
												localparam VX_gpu_pkg_EX_TCU = 2;
												localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
												localparam VX_gpu_pkg_EX_BITS = 2;
												localparam VX_gpu_pkg_INST_OP_BITS = 4;
												localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
												localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
												localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_RV_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
												localparam VX_gpu_pkg_PC_BITS = 30;
												localparam VX_gpu_pkg_SIMD_COUNT = 1;
												localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
												localparam VX_gpu_pkg_SIMD_IDX_W = 1;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
												// removed localparam type VX_gpu_pkg_alu_args_t
												localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
												// removed localparam type VX_gpu_pkg_csr_args_t
												localparam VX_gpu_pkg_INST_FMT_BITS = 2;
												localparam VX_gpu_pkg_INST_FRM_BITS = 3;
												// removed localparam type VX_gpu_pkg_fpu_args_t
												localparam VX_gpu_pkg_OFFSET_BITS = 12;
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												// removed localparam type VX_gpu_pkg_operands_t
												wire [472:0] data;
												// Trace: src/VX_operands_if.sv:4:5
												wire ready;
												// Trace: src/VX_operands_if.sv:5:5
												// Trace: src/VX_operands_if.sv:10:5
											end
											// Trace: src/VX_issue_slice.sv:15:5
											// expanded module instance: ibuffer
											localparam _bbase_D579A_ibuffer_if = 0;
											localparam _param_D579A_INSTANCE_ID = "";
											localparam _param_D579A_ISSUE_ID = ISSUE_ID;
											if (1) begin : ibuffer
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_ibuffer.sv:2:15
												localparam INSTANCE_ID = _param_D579A_INSTANCE_ID;
												// Trace: src/VX_ibuffer.sv:3:15
												localparam ISSUE_ID = _param_D579A_ISSUE_ID;
												// Trace: src/VX_ibuffer.sv:5:5
												wire clk;
												// Trace: src/VX_ibuffer.sv:6:5
												wire reset;
												// Trace: src/VX_ibuffer.sv:7:5
												// removed modport instance decode_if
												// Trace: src/VX_ibuffer.sv:8:5
												localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
												localparam _mbase_ibuffer_if = 0;
												// Trace: src/VX_ibuffer.sv:10:5
												localparam VX_gpu_pkg_EX_SFU = 2;
												localparam VX_gpu_pkg_EX_FPU = 2;
												localparam VX_gpu_pkg_EX_TCU = 2;
												localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
												localparam VX_gpu_pkg_EX_BITS = 2;
												localparam VX_gpu_pkg_INST_OP_BITS = 4;
												localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
												localparam VX_gpu_pkg_PC_BITS = 30;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
												// removed localparam type VX_gpu_pkg_alu_args_t
												localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
												// removed localparam type VX_gpu_pkg_csr_args_t
												localparam VX_gpu_pkg_INST_FMT_BITS = 2;
												localparam VX_gpu_pkg_INST_FRM_BITS = 3;
												// removed localparam type VX_gpu_pkg_fpu_args_t
												localparam VX_gpu_pkg_OFFSET_BITS = 12;
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_REG_TYPE_BITS = 1;
												localparam VX_gpu_pkg_RV_REGS_BITS = 5;
												// removed localparam type VX_gpu_pkg_reg_idx_t
												// removed localparam type VX_gpu_pkg_ibuffer_t
												localparam OUT_DATAW = 106;
												// Trace: src/VX_ibuffer.sv:11:5
												localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
												localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
												localparam VX_gpu_pkg_ISSUE_ISW_BITS = 0;
												localparam VX_gpu_pkg_NW_BITS = 2;
												localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
												function automatic [1:0] VX_gpu_pkg_wid_to_wis;
													// Trace: src/VX_gpu_pkg.sv:285:9
													input reg [1:0] wid;
													// Trace: src/VX_gpu_pkg.sv:287:9
													begin
														// Trace: src/VX_gpu_pkg.sv:288:13
														VX_gpu_pkg_wid_to_wis = wid >> VX_gpu_pkg_ISSUE_ISW_BITS;
													end
												endfunction
												wire [1:0] decode_wis = VX_gpu_pkg_wid_to_wis(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[106-:2]);
												// Trace: src/VX_ibuffer.sv:12:5
												wire [3:0] ibuf_ready_in;
												// Trace: src/VX_ibuffer.sv:13:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.ready = ibuf_ready_in[decode_wis];
												// Trace: src/VX_ibuffer.sv:14:5
												genvar _gv_w_1;
												for (_gv_w_1 = 0; _gv_w_1 < VX_gpu_pkg_PER_ISSUE_WARPS; _gv_w_1 = _gv_w_1 + 1) begin : g_instr_bufs
													localparam w = _gv_w_1;
													// Trace: src/VX_ibuffer.sv:15:9
													// expanded interface instance: uop_sequencer_if
													if (1) begin : uop_sequencer_if
														// removed import VX_gpu_pkg::*;
														// Trace: src/VX_ibuffer_if.sv:2:5
														wire valid;
														// Trace: src/VX_ibuffer_if.sv:3:5
														localparam VX_gpu_pkg_EX_SFU = 2;
														localparam VX_gpu_pkg_EX_FPU = 2;
														localparam VX_gpu_pkg_EX_TCU = 2;
														localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
														localparam VX_gpu_pkg_EX_BITS = 2;
														localparam VX_gpu_pkg_INST_OP_BITS = 4;
														localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
														localparam VX_gpu_pkg_PC_BITS = 30;
														localparam VX_gpu_pkg_UUID_WIDTH = 1;
														localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
														// removed localparam type VX_gpu_pkg_alu_args_t
														localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
														// removed localparam type VX_gpu_pkg_csr_args_t
														localparam VX_gpu_pkg_INST_FMT_BITS = 2;
														localparam VX_gpu_pkg_INST_FRM_BITS = 3;
														// removed localparam type VX_gpu_pkg_fpu_args_t
														localparam VX_gpu_pkg_OFFSET_BITS = 12;
														// removed localparam type VX_gpu_pkg_lsu_args_t
														// removed localparam type VX_gpu_pkg_wctl_args_t
														// removed localparam type VX_gpu_pkg_op_args_t
														localparam VX_gpu_pkg_REG_TYPES = 1;
														localparam VX_gpu_pkg_REG_TYPE_BITS = 1;
														localparam VX_gpu_pkg_RV_REGS_BITS = 5;
														// removed localparam type VX_gpu_pkg_reg_idx_t
														// removed localparam type VX_gpu_pkg_ibuffer_t
														wire [105:0] data;
														// Trace: src/VX_ibuffer_if.sv:4:5
														wire ready;
														// Trace: src/VX_ibuffer_if.sv:5:5
														// Trace: src/VX_ibuffer_if.sv:10:5
													end
													// Trace: src/VX_ibuffer.sv:16:9
													VX_elastic_buffer #(
														.DATAW(OUT_DATAW),
														.SIZE(4),
														.OUT_REG(1)
													) instr_buf(
														.clk(clk),
														.reset(reset),
														.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.valid && (decode_wis == sv2v_cast_2_signed(w))),
														.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[107], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[104-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[100-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[70-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[68-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[64-:37], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[27], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[26-:3], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[23-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[17-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[11-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].slice_decode_if.data[5-:6]}),
														.ready_in(ibuf_ready_in[w]),
														.valid_out(uop_sequencer_if.valid),
														.data_out(uop_sequencer_if.data),
														.ready_out(uop_sequencer_if.ready)
													);
													// Trace: src/VX_ibuffer.sv:43:9
													// expanded module instance: uop_sequencer
													localparam _bbase_70C82_output_if = w + _mbase_ibuffer_if;
													if (1) begin : uop_sequencer
														// removed import VX_gpu_pkg::*;
														// Trace: src/VX_uop_sequencer.sv:3:5
														wire clk;
														// Trace: src/VX_uop_sequencer.sv:4:5
														wire reset;
														// Trace: src/VX_uop_sequencer.sv:5:5
														// removed modport instance input_if
														// Trace: src/VX_uop_sequencer.sv:6:5
														localparam _mbase_output_if = _bbase_70C82_output_if;
														// Trace: src/VX_uop_sequencer.sv:8:5
														localparam VX_gpu_pkg_EX_SFU = 2;
														localparam VX_gpu_pkg_EX_FPU = 2;
														localparam VX_gpu_pkg_EX_TCU = 2;
														localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
														localparam VX_gpu_pkg_EX_BITS = 2;
														localparam VX_gpu_pkg_INST_OP_BITS = 4;
														localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
														localparam VX_gpu_pkg_PC_BITS = 30;
														localparam VX_gpu_pkg_UUID_WIDTH = 1;
														localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
														// removed localparam type VX_gpu_pkg_alu_args_t
														localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
														// removed localparam type VX_gpu_pkg_csr_args_t
														localparam VX_gpu_pkg_INST_FMT_BITS = 2;
														localparam VX_gpu_pkg_INST_FRM_BITS = 3;
														// removed localparam type VX_gpu_pkg_fpu_args_t
														localparam VX_gpu_pkg_OFFSET_BITS = 12;
														// removed localparam type VX_gpu_pkg_lsu_args_t
														// removed localparam type VX_gpu_pkg_wctl_args_t
														// removed localparam type VX_gpu_pkg_op_args_t
														localparam VX_gpu_pkg_REG_TYPES = 1;
														localparam VX_gpu_pkg_REG_TYPE_BITS = 1;
														localparam VX_gpu_pkg_RV_REGS_BITS = 5;
														// removed localparam type VX_gpu_pkg_reg_idx_t
														// removed localparam type VX_gpu_pkg_ibuffer_t
														wire [105:0] uop_data;
														// Trace: src/VX_uop_sequencer.sv:9:5
														wire is_uop_input;
														// Trace: src/VX_uop_sequencer.sv:10:5
														wire uop_start = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer.g_instr_bufs[_gv_w_1].uop_sequencer_if.valid && is_uop_input;
														// Trace: src/VX_uop_sequencer.sv:11:5
														wire uop_next = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[_mbase_output_if].ready;
														// Trace: src/VX_uop_sequencer.sv:12:5
														wire uop_done;
														// Trace: src/VX_uop_sequencer.sv:13:5
														assign is_uop_input = 0;
														// Trace: src/VX_uop_sequencer.sv:14:5
														assign uop_done = 0;
														// Trace: src/VX_uop_sequencer.sv:15:5
														assign uop_data = 1'sb0;
														// Trace: src/VX_uop_sequencer.sv:16:5
														reg uop_active;
														// Trace: src/VX_uop_sequencer.sv:17:5
														always @(posedge clk)
															// Trace: src/VX_uop_sequencer.sv:18:9
															if (reset)
																// Trace: src/VX_uop_sequencer.sv:19:13
																uop_active <= 0;
															else
																// Trace: src/VX_uop_sequencer.sv:21:13
																if (uop_active) begin
																	begin
																		// Trace: src/VX_uop_sequencer.sv:22:17
																		if (uop_next && uop_done)
																			// Trace: src/VX_uop_sequencer.sv:23:21
																			uop_active <= 0;
																	end
																end
																else if (uop_start)
																	// Trace: src/VX_uop_sequencer.sv:27:17
																	uop_active <= 1;
														// Trace: src/VX_uop_sequencer.sv:31:5
														wire uop_hold = ~uop_active && is_uop_input;
														// Trace: src/VX_uop_sequencer.sv:32:5
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[_mbase_output_if].valid = (uop_active ? 1'b1 : Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer.g_instr_bufs[_gv_w_1].uop_sequencer_if.valid && ~uop_hold);
														// Trace: src/VX_uop_sequencer.sv:33:5
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[_mbase_output_if].data = (uop_active ? uop_data : Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer.g_instr_bufs[_gv_w_1].uop_sequencer_if.data);
														// Trace: src/VX_uop_sequencer.sv:34:5
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer.g_instr_bufs[_gv_w_1].uop_sequencer_if.ready = (uop_active ? Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[_mbase_output_if].ready && uop_done : Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[_mbase_output_if].ready && ~uop_hold);
													end
													assign uop_sequencer.clk = clk;
													assign uop_sequencer.reset = reset;
												end
											end
											assign ibuffer.clk = clk;
											assign ibuffer.reset = reset;
											// Trace: src/VX_issue_slice.sv:24:5
											// expanded module instance: scoreboard
											localparam _bbase_85D2C_writeback_if = issue_id + _mbase_writeback_if;
											localparam _bbase_85D2C_ibuffer_if = 0;
											localparam _param_85D2C_INSTANCE_ID = "";
											localparam _param_85D2C_ISSUE_ID = ISSUE_ID;
											if (1) begin : scoreboard
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_scoreboard.sv:2:15
												localparam INSTANCE_ID = _param_85D2C_INSTANCE_ID;
												// Trace: src/VX_scoreboard.sv:3:15
												localparam ISSUE_ID = _param_85D2C_ISSUE_ID;
												// Trace: src/VX_scoreboard.sv:5:5
												wire clk;
												// Trace: src/VX_scoreboard.sv:6:5
												wire reset;
												// Trace: src/VX_scoreboard.sv:7:5
												localparam _mbase_writeback_if = _bbase_85D2C_writeback_if;
												// Trace: src/VX_scoreboard.sv:8:5
												localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
												localparam _mbase_ibuffer_if = 0;
												// Trace: src/VX_scoreboard.sv:9:5
												// removed modport instance scoreboard_if
												// Trace: src/VX_scoreboard.sv:11:5
												localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
												localparam NUM_OPDS = 4;
												// Trace: src/VX_scoreboard.sv:12:5
												localparam VX_gpu_pkg_EX_SFU = 2;
												localparam VX_gpu_pkg_EX_FPU = 2;
												localparam VX_gpu_pkg_EX_TCU = 2;
												localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
												localparam VX_gpu_pkg_EX_BITS = 2;
												localparam VX_gpu_pkg_INST_OP_BITS = 4;
												localparam VX_gpu_pkg_PC_BITS = 30;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
												// removed localparam type VX_gpu_pkg_alu_args_t
												localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
												// removed localparam type VX_gpu_pkg_csr_args_t
												localparam VX_gpu_pkg_INST_FMT_BITS = 2;
												localparam VX_gpu_pkg_INST_FRM_BITS = 3;
												// removed localparam type VX_gpu_pkg_fpu_args_t
												localparam VX_gpu_pkg_OFFSET_BITS = 12;
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_REG_TYPE_BITS = 1;
												localparam VX_gpu_pkg_RV_REGS_BITS = 5;
												// removed localparam type VX_gpu_pkg_reg_idx_t
												// removed localparam type VX_gpu_pkg_ibuffer_t
												localparam IN_DATAW = 106;
												// Trace: src/VX_scoreboard.sv:13:5
												// expanded interface instance: staging_if
												genvar _arr_8EA22;
												for (_arr_8EA22 = 0; _arr_8EA22 <= 3; _arr_8EA22 = _arr_8EA22 + 1) begin : staging_if
													// removed import VX_gpu_pkg::*;
													// Trace: src/VX_ibuffer_if.sv:2:5
													wire valid;
													// Trace: src/VX_ibuffer_if.sv:3:5
													localparam VX_gpu_pkg_EX_SFU = 2;
													localparam VX_gpu_pkg_EX_FPU = 2;
													localparam VX_gpu_pkg_EX_TCU = 2;
													localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
													localparam VX_gpu_pkg_EX_BITS = 2;
													localparam VX_gpu_pkg_INST_OP_BITS = 4;
													localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
													localparam VX_gpu_pkg_PC_BITS = 30;
													localparam VX_gpu_pkg_UUID_WIDTH = 1;
													localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
													// removed localparam type VX_gpu_pkg_alu_args_t
													localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
													// removed localparam type VX_gpu_pkg_csr_args_t
													localparam VX_gpu_pkg_INST_FMT_BITS = 2;
													localparam VX_gpu_pkg_INST_FRM_BITS = 3;
													// removed localparam type VX_gpu_pkg_fpu_args_t
													localparam VX_gpu_pkg_OFFSET_BITS = 12;
													// removed localparam type VX_gpu_pkg_lsu_args_t
													// removed localparam type VX_gpu_pkg_wctl_args_t
													// removed localparam type VX_gpu_pkg_op_args_t
													localparam VX_gpu_pkg_REG_TYPES = 1;
													localparam VX_gpu_pkg_REG_TYPE_BITS = 1;
													localparam VX_gpu_pkg_RV_REGS_BITS = 5;
													// removed localparam type VX_gpu_pkg_reg_idx_t
													// removed localparam type VX_gpu_pkg_ibuffer_t
													wire [105:0] data;
													// Trace: src/VX_ibuffer_if.sv:4:5
													wire ready;
													// Trace: src/VX_ibuffer_if.sv:5:5
													// Trace: src/VX_ibuffer_if.sv:10:5
												end
												// Trace: src/VX_scoreboard.sv:14:5
												wire [3:0] operands_ready;
												// Trace: src/VX_scoreboard.sv:15:5
												genvar _gv_w_2;
												for (_gv_w_2 = 0; _gv_w_2 < VX_gpu_pkg_PER_ISSUE_WARPS; _gv_w_2 = _gv_w_2 + 1) begin : g_stanging_bufs
													localparam w = _gv_w_2;
													// Trace: src/VX_scoreboard.sv:16:9
													VX_pipe_buffer #(.DATAW(IN_DATAW)) stanging_buf(
														.clk(clk),
														.reset(reset),
														.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].valid),
														.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data),
														.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].ready),
														.valid_out(staging_if[w].valid),
														.data_out(staging_if[w].data),
														.ready_out(staging_if[w].ready)
													);
												end
												// Trace: src/VX_scoreboard.sv:29:5
												genvar _gv_w_3;
												localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
												localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
												localparam VX_gpu_pkg_RV_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS = 32;
												function automatic [31:0] VX_gpu_pkg_to_reg_mask;
													// Trace: src/VX_gpu_pkg.sv:595:56
													input reg [5:0] reg_idx;
													// Trace: src/VX_gpu_pkg.sv:596:9
													VX_gpu_pkg_to_reg_mask = 1 << reg_idx[4-:5];
												endfunction
												for (_gv_w_3 = 0; _gv_w_3 < VX_gpu_pkg_PER_ISSUE_WARPS; _gv_w_3 = _gv_w_3 + 1) begin : g_scoreboard
													localparam w = _gv_w_3;
													// Trace: src/VX_scoreboard.sv:30:9
													reg [31:0] inuse_regs;
													reg [31:0] inuse_regs_n;
													// Trace: src/VX_scoreboard.sv:31:9
													wire [3:0] operands_busy;
													// Trace: src/VX_scoreboard.sv:32:9
													wire ibuffer_fire = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].ready;
													// Trace: src/VX_scoreboard.sv:33:9
													wire staging_fire = staging_if[w].valid && staging_if[w].ready;
													// Trace: src/VX_scoreboard.sv:34:9
													wire writeback_fire = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].valid && (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[171-:2] == sv2v_cast_2_signed(w))) && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[0];
													// Trace: src/VX_scoreboard.sv:37:9
													wire [23:0] ibf_opds;
													wire [23:0] stg_opds;
													// Trace: src/VX_scoreboard.sv:38:9
													assign ibf_opds = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data[5-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data[11-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data[17-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data[23-:6]};
													// Trace: src/VX_scoreboard.sv:39:9
													assign stg_opds = {staging_if[w].data[5-:6], staging_if[w].data[11-:6], staging_if[w].data[17-:6], staging_if[w].data[23-:6]};
													// Trace: src/VX_scoreboard.sv:40:9
													wire [3:0] ibf_used_rs = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data[26-:3], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.ibuffer_if[w + _mbase_ibuffer_if].data[27]};
													// Trace: src/VX_scoreboard.sv:41:9
													wire [3:0] stg_used_rs = {staging_if[w].data[26-:3], staging_if[w].data[27]};
													// Trace: src/VX_scoreboard.sv:42:9
													wire [127:0] ibf_opd_mask;
													wire [127:0] stg_opd_mask;
													genvar _gv_i_134;
													for (_gv_i_134 = 0; _gv_i_134 < NUM_OPDS; _gv_i_134 = _gv_i_134 + 1) begin : g_opd_masks
														localparam i = _gv_i_134;
														genvar _gv_j_16;
														for (_gv_j_16 = 0; _gv_j_16 < VX_gpu_pkg_REG_TYPES; _gv_j_16 = _gv_j_16 + 1) begin : g_j
															localparam j = _gv_j_16;
															// Trace: src/VX_scoreboard.sv:45:17
															assign ibf_opd_mask[(i + j) * 32+:32] = VX_gpu_pkg_to_reg_mask(ibf_opds[i * 6+:6]) & {VX_gpu_pkg_RV_REGS {ibf_used_rs[i] && (ibf_opds[(i * 6) + 5-:1] == j)}};
															// Trace: src/VX_scoreboard.sv:46:17
															assign stg_opd_mask[(i + j) * 32+:32] = VX_gpu_pkg_to_reg_mask(stg_opds[i * 6+:6]) & {VX_gpu_pkg_RV_REGS {stg_used_rs[i] && (stg_opds[(i * 6) + 5-:1] == j)}};
														end
													end
													// Trace: src/VX_scoreboard.sv:49:9
													always @(*) begin
														// Trace: src/VX_scoreboard.sv:50:13
														inuse_regs_n = inuse_regs;
														// Trace: src/VX_scoreboard.sv:51:13
														if (writeback_fire)
															// Trace: src/VX_scoreboard.sv:52:17
															inuse_regs_n[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data[134-:5]] = 0;
														if (staging_fire && staging_if[w].data[27])
															// Trace: src/VX_scoreboard.sv:55:17
															inuse_regs_n = inuse_regs_n | stg_opd_mask[0+:32];
													end
													// Trace: src/VX_scoreboard.sv:58:9
													wire [31:0] in_use_mask;
													genvar _gv_i_135;
													for (_gv_i_135 = 0; _gv_i_135 < VX_gpu_pkg_REG_TYPES; _gv_i_135 = _gv_i_135 + 1) begin : g_in_use_mask
														localparam i = _gv_i_135;
														// Trace: src/VX_scoreboard.sv:60:13
														wire [31:0] ibf_reg_mask = ((ibf_opd_mask[i * 32+:32] | ibf_opd_mask[(1 + i) * 32+:32]) | ibf_opd_mask[(2 + i) * 32+:32]) | ibf_opd_mask[(3 + i) * 32+:32];
														// Trace: src/VX_scoreboard.sv:61:13
														wire [31:0] stg_reg_mask = ((stg_opd_mask[i * 32+:32] | stg_opd_mask[(1 + i) * 32+:32]) | stg_opd_mask[(2 + i) * 32+:32]) | stg_opd_mask[(3 + i) * 32+:32];
														// Trace: src/VX_scoreboard.sv:62:13
														wire [31:0] regs_mask = (ibuffer_fire ? ibf_reg_mask : stg_reg_mask);
														// Trace: src/VX_scoreboard.sv:63:13
														assign in_use_mask[i * 32+:32] = inuse_regs_n[i * VX_gpu_pkg_RV_REGS+:VX_gpu_pkg_RV_REGS] & regs_mask;
													end
													// Trace: src/VX_scoreboard.sv:65:9
													wire [0:0] regs_busy;
													genvar _gv_i_136;
													for (_gv_i_136 = 0; _gv_i_136 < VX_gpu_pkg_REG_TYPES; _gv_i_136 = _gv_i_136 + 1) begin : g_regs_busy
														localparam i = _gv_i_136;
														// Trace: src/VX_scoreboard.sv:67:13
														assign regs_busy[i] = in_use_mask[i * 32+:32] != 0;
													end
													genvar _gv_i_137;
													for (_gv_i_137 = 0; _gv_i_137 < NUM_OPDS; _gv_i_137 = _gv_i_137 + 1) begin : g_operands_busy
														localparam i = _gv_i_137;
														// Trace: src/VX_scoreboard.sv:70:13
														wire [0:0] rtype = stg_opds[(i * 6) + 5-:1];
														// Trace: src/VX_scoreboard.sv:71:13
														assign operands_busy[i] = (in_use_mask[rtype * 32+:32] & stg_opd_mask[(i + rtype) * 32+:32]) != 0;
													end
													// Trace: src/VX_scoreboard.sv:73:9
													reg operands_ready_r;
													// Trace: src/VX_scoreboard.sv:74:9
													always @(posedge clk) begin
														// Trace: src/VX_scoreboard.sv:75:13
														if (reset)
															// Trace: src/VX_scoreboard.sv:76:17
															inuse_regs <= 1'sb0;
														else
															// Trace: src/VX_scoreboard.sv:78:17
															inuse_regs <= inuse_regs_n;
														// Trace: src/VX_scoreboard.sv:80:13
														operands_ready_r <= ~(|regs_busy);
													end
													// Trace: src/VX_scoreboard.sv:82:9
													assign operands_ready[w] = operands_ready_r;
												end
												// Trace: src/VX_scoreboard.sv:84:5
												wire [3:0] arb_valid_in;
												// Trace: src/VX_scoreboard.sv:85:5
												wire [423:0] arb_data_in;
												// Trace: src/VX_scoreboard.sv:86:5
												wire [3:0] arb_ready_in;
												// Trace: src/VX_scoreboard.sv:87:5
												genvar _gv_w_4;
												for (_gv_w_4 = 0; _gv_w_4 < VX_gpu_pkg_PER_ISSUE_WARPS; _gv_w_4 = _gv_w_4 + 1) begin : g_arb_data_in
													localparam w = _gv_w_4;
													// Trace: src/VX_scoreboard.sv:88:9
													assign arb_valid_in[w] = staging_if[w].valid && operands_ready[w];
													// Trace: src/VX_scoreboard.sv:89:9
													assign arb_data_in[w * 106+:106] = staging_if[w].data;
													// Trace: src/VX_scoreboard.sv:90:9
													assign staging_if[w].ready = arb_ready_in[w] && operands_ready[w];
												end
												// Trace: src/VX_scoreboard.sv:92:5
												VX_stream_arb #(
													.NUM_INPUTS(VX_gpu_pkg_PER_ISSUE_WARPS),
													.DATAW(IN_DATAW),
													.ARBITER("C"),
													.OUT_BUF(3)
												) out_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(arb_valid_in),
													.ready_in(arb_ready_in),
													.data_in(arb_data_in),
													.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[107], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[104-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[100-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[70-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[68-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[64-:37], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[27], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[26-:3], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[23-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[17-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[11-:6], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[5-:6]}),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.ready),
													.sel_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data[106-:2])
												);
											end
											assign scoreboard.clk = clk;
											assign scoreboard.reset = reset;
											// Trace: src/VX_issue_slice.sv:34:5
											// expanded module instance: operands
											localparam _bbase_CD6E0_writeback_if = issue_id + _mbase_writeback_if;
											localparam _param_CD6E0_INSTANCE_ID = "";
											localparam _param_CD6E0_ISSUE_ID = ISSUE_ID;
											if (1) begin : operands
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_operands.sv:2:15
												localparam INSTANCE_ID = _param_CD6E0_INSTANCE_ID;
												// Trace: src/VX_operands.sv:3:15
												localparam ISSUE_ID = _param_CD6E0_ISSUE_ID;
												// Trace: src/VX_operands.sv:5:5
												wire clk;
												// Trace: src/VX_operands.sv:6:5
												wire reset;
												// Trace: src/VX_operands.sv:7:5
												localparam _mbase_writeback_if = _bbase_CD6E0_writeback_if;
												// Trace: src/VX_operands.sv:8:5
												// removed modport instance scoreboard_if
												// Trace: src/VX_operands.sv:9:5
												// removed modport instance operands_if
												// Trace: src/VX_operands.sv:11:5
												localparam VX_gpu_pkg_EX_SFU = 2;
												localparam VX_gpu_pkg_EX_FPU = 2;
												localparam VX_gpu_pkg_EX_TCU = 2;
												localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
												localparam VX_gpu_pkg_EX_BITS = 2;
												localparam VX_gpu_pkg_INST_OP_BITS = 4;
												localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
												localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
												localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_RV_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
												localparam VX_gpu_pkg_PC_BITS = 30;
												localparam VX_gpu_pkg_SIMD_COUNT = 1;
												localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
												localparam VX_gpu_pkg_SIMD_IDX_W = 1;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
												// removed localparam type VX_gpu_pkg_alu_args_t
												localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
												// removed localparam type VX_gpu_pkg_csr_args_t
												localparam VX_gpu_pkg_INST_FMT_BITS = 2;
												localparam VX_gpu_pkg_INST_FRM_BITS = 3;
												// removed localparam type VX_gpu_pkg_fpu_args_t
												localparam VX_gpu_pkg_OFFSET_BITS = 12;
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												// removed localparam type VX_gpu_pkg_operands_t
												localparam OUT_DATAW = 473;
												// Trace: src/VX_operands.sv:12:5
												localparam OUT_ARB_STICKY = 1'd0;
												// Trace: src/VX_operands.sv:13:5
												// expanded interface instance: per_opc_operands_if
												genvar _arr_C37C1;
												for (_arr_C37C1 = 0; _arr_C37C1 <= 0; _arr_C37C1 = _arr_C37C1 + 1) begin : per_opc_operands_if
													// removed import VX_gpu_pkg::*;
													// Trace: src/VX_operands_if.sv:2:5
													wire valid;
													// Trace: src/VX_operands_if.sv:3:5
													localparam VX_gpu_pkg_EX_SFU = 2;
													localparam VX_gpu_pkg_EX_FPU = 2;
													localparam VX_gpu_pkg_EX_TCU = 2;
													localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
													localparam VX_gpu_pkg_EX_BITS = 2;
													localparam VX_gpu_pkg_INST_OP_BITS = 4;
													localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
													localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
													localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
													localparam VX_gpu_pkg_REG_TYPES = 1;
													localparam VX_gpu_pkg_RV_REGS = 32;
													localparam VX_gpu_pkg_NUM_REGS = 32;
													localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
													localparam VX_gpu_pkg_PC_BITS = 30;
													localparam VX_gpu_pkg_SIMD_COUNT = 1;
													localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
													localparam VX_gpu_pkg_SIMD_IDX_W = 1;
													localparam VX_gpu_pkg_UUID_WIDTH = 1;
													localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
													// removed localparam type VX_gpu_pkg_alu_args_t
													localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
													// removed localparam type VX_gpu_pkg_csr_args_t
													localparam VX_gpu_pkg_INST_FMT_BITS = 2;
													localparam VX_gpu_pkg_INST_FRM_BITS = 3;
													// removed localparam type VX_gpu_pkg_fpu_args_t
													localparam VX_gpu_pkg_OFFSET_BITS = 12;
													// removed localparam type VX_gpu_pkg_lsu_args_t
													// removed localparam type VX_gpu_pkg_wctl_args_t
													// removed localparam type VX_gpu_pkg_op_args_t
													// removed localparam type VX_gpu_pkg_operands_t
													wire [472:0] data;
													// Trace: src/VX_operands_if.sv:4:5
													wire ready;
													// Trace: src/VX_operands_if.sv:5:5
													// Trace: src/VX_operands_if.sv:10:5
												end
												// Trace: src/VX_operands.sv:14:5
												localparam VX_gpu_pkg_NUM_OPCS_BITS = 0;
												localparam VX_gpu_pkg_NUM_OPCS_W = 1;
												wire [0:0] sb_opc;
												wire [0:0] wb_opc;
												// Trace: src/VX_operands.sv:15:5
												if (1) begin : g_wis_opc
													// Trace: src/VX_operands.sv:19:9
													assign sb_opc = 0;
													// Trace: src/VX_operands.sv:20:9
													assign wb_opc = 0;
												end
												// Trace: src/VX_operands.sv:22:5
												wire [0:0] scoreboard_ready_in;
												// Trace: src/VX_operands.sv:23:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.ready = scoreboard_ready_in[sb_opc];
												// Trace: src/VX_operands.sv:24:5
												genvar _gv_i_206;
												for (_gv_i_206 = 0; _gv_i_206 < 1; _gv_i_206 = _gv_i_206 + 1) begin : g_collectors
													localparam i = _gv_i_206;
													// Trace: src/VX_operands.sv:25:9
													// expanded interface instance: opc_scoreboard_if
													if (1) begin : opc_scoreboard_if
														// removed import VX_gpu_pkg::*;
														// Trace: src/VX_scoreboard_if.sv:2:5
														wire valid;
														// Trace: src/VX_scoreboard_if.sv:3:5
														localparam VX_gpu_pkg_EX_SFU = 2;
														localparam VX_gpu_pkg_EX_FPU = 2;
														localparam VX_gpu_pkg_EX_TCU = 2;
														localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
														localparam VX_gpu_pkg_EX_BITS = 2;
														localparam VX_gpu_pkg_INST_OP_BITS = 4;
														localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
														localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
														localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
														localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
														localparam VX_gpu_pkg_PC_BITS = 30;
														localparam VX_gpu_pkg_UUID_WIDTH = 1;
														localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
														// removed localparam type VX_gpu_pkg_alu_args_t
														localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
														// removed localparam type VX_gpu_pkg_csr_args_t
														localparam VX_gpu_pkg_INST_FMT_BITS = 2;
														localparam VX_gpu_pkg_INST_FRM_BITS = 3;
														// removed localparam type VX_gpu_pkg_fpu_args_t
														localparam VX_gpu_pkg_OFFSET_BITS = 12;
														// removed localparam type VX_gpu_pkg_lsu_args_t
														// removed localparam type VX_gpu_pkg_wctl_args_t
														// removed localparam type VX_gpu_pkg_op_args_t
														localparam VX_gpu_pkg_REG_TYPES = 1;
														localparam VX_gpu_pkg_REG_TYPE_BITS = 1;
														localparam VX_gpu_pkg_RV_REGS_BITS = 5;
														// removed localparam type VX_gpu_pkg_reg_idx_t
														// removed localparam type VX_gpu_pkg_scoreboard_t
														wire [107:0] data;
														// Trace: src/VX_scoreboard_if.sv:4:5
														wire ready;
														// Trace: src/VX_scoreboard_if.sv:5:5
														// Trace: src/VX_scoreboard_if.sv:10:5
													end
													// Trace: src/VX_operands.sv:26:9
													assign opc_scoreboard_if.valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.valid && (sb_opc == i);
													// Trace: src/VX_operands.sv:27:9
													assign opc_scoreboard_if.data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.scoreboard_if.data;
													// Trace: src/VX_operands.sv:28:9
													assign scoreboard_ready_in[i] = opc_scoreboard_if.ready;
													// Trace: src/VX_operands.sv:29:9
													// expanded interface instance: opc_writeback_if
													if (1) begin : opc_writeback_if
														// removed import VX_gpu_pkg::*;
														// Trace: src/VX_writeback_if.sv:2:5
														wire valid;
														// Trace: src/VX_writeback_if.sv:3:5
														localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
														localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
														localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
														localparam VX_gpu_pkg_REG_TYPES = 1;
														localparam VX_gpu_pkg_RV_REGS = 32;
														localparam VX_gpu_pkg_NUM_REGS = 32;
														localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
														localparam VX_gpu_pkg_PC_BITS = 30;
														localparam VX_gpu_pkg_SIMD_COUNT = 1;
														localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
														localparam VX_gpu_pkg_SIMD_IDX_W = 1;
														localparam VX_gpu_pkg_UUID_WIDTH = 1;
														// removed localparam type VX_gpu_pkg_writeback_t
														wire [172:0] data;
														// Trace: src/VX_writeback_if.sv:4:5
														// Trace: src/VX_writeback_if.sv:8:5
													end
													// Trace: src/VX_operands.sv:30:9
													assign opc_writeback_if.valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].valid && (wb_opc == i);
													// Trace: src/VX_operands.sv:31:9
													assign opc_writeback_if.data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[_mbase_writeback_if].data;
													// Trace: src/VX_operands.sv:32:9
													// expanded module instance: opc_unit
													localparam _bbase_A91FA_operands_if = i;
													localparam _param_A91FA_INSTANCE_ID = "";
													localparam _param_A91FA_NUM_BANKS = 4;
													localparam _param_A91FA_OUT_BUF = 3;
													if (1) begin : opc_unit
														// removed import VX_gpu_pkg::*;
														// Trace: src/VX_opc_unit.sv:2:15
														localparam INSTANCE_ID = _param_A91FA_INSTANCE_ID;
														// Trace: src/VX_opc_unit.sv:3:15
														localparam NUM_BANKS = _param_A91FA_NUM_BANKS;
														// Trace: src/VX_opc_unit.sv:4:15
														localparam OUT_BUF = _param_A91FA_OUT_BUF;
														// Trace: src/VX_opc_unit.sv:6:5
														wire clk;
														// Trace: src/VX_opc_unit.sv:7:5
														wire reset;
														// Trace: src/VX_opc_unit.sv:8:5
														// removed modport instance writeback_if
														// Trace: src/VX_opc_unit.sv:9:5
														// removed modport instance scoreboard_if
														// Trace: src/VX_opc_unit.sv:10:5
														localparam _mbase_operands_if = _bbase_A91FA_operands_if;
														// Trace: src/VX_opc_unit.sv:12:5
														localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
														localparam VX_gpu_pkg_SRC_OPD_BITS = 2;
														localparam VX_gpu_pkg_SRC_OPD_WIDTH = VX_gpu_pkg_SRC_OPD_BITS;
														localparam REQ_SEL_WIDTH = VX_gpu_pkg_SRC_OPD_WIDTH;
														// Trace: src/VX_opc_unit.sv:13:5
														localparam BANK_SEL_BITS = 2;
														// Trace: src/VX_opc_unit.sv:14:5
														localparam BANK_SEL_WIDTH = BANK_SEL_BITS;
														// Trace: src/VX_opc_unit.sv:15:5
														localparam BANK_DATA_WIDTH = 128;
														// Trace: src/VX_opc_unit.sv:16:5
														localparam BANK_DATA_SIZE = 16;
														// Trace: src/VX_opc_unit.sv:17:5
														localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
														localparam PER_OPC_WARPS = 4;
														// Trace: src/VX_opc_unit.sv:18:5
														localparam PER_OPC_NW_BITS = 2;
														// Trace: src/VX_opc_unit.sv:19:5
														localparam VX_gpu_pkg_REG_TYPES = 1;
														localparam VX_gpu_pkg_RV_REGS = 32;
														localparam VX_gpu_pkg_NUM_REGS = 32;
														localparam VX_gpu_pkg_SIMD_COUNT = 1;
														localparam BANK_SIZE = 32;
														// Trace: src/VX_opc_unit.sv:20:5
														localparam BANK_ADDR_WIDTH = 5;
														// Trace: src/VX_opc_unit.sv:21:5
														localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
														localparam REG_REM_BITS = 3;
														// Trace: src/VX_opc_unit.sv:22:5
														localparam VX_gpu_pkg_EX_SFU = 2;
														localparam VX_gpu_pkg_EX_FPU = 2;
														localparam VX_gpu_pkg_EX_TCU = 2;
														localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
														localparam VX_gpu_pkg_EX_BITS = 2;
														localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
														localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
														localparam VX_gpu_pkg_INST_OP_BITS = 4;
														localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
														localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
														localparam VX_gpu_pkg_PC_BITS = 30;
														localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
														localparam VX_gpu_pkg_SIMD_IDX_W = 1;
														localparam VX_gpu_pkg_UUID_WIDTH = 1;
														localparam META_DATAW = 89;
														// Trace: src/VX_opc_unit.sv:23:5
														// removed localparam type VX_gpu_pkg_alu_args_t
														// removed localparam type VX_gpu_pkg_csr_args_t
														localparam VX_gpu_pkg_INST_FMT_BITS = 2;
														localparam VX_gpu_pkg_INST_FRM_BITS = 3;
														// removed localparam type VX_gpu_pkg_fpu_args_t
														localparam VX_gpu_pkg_OFFSET_BITS = 12;
														// removed localparam type VX_gpu_pkg_lsu_args_t
														// removed localparam type VX_gpu_pkg_wctl_args_t
														// removed localparam type VX_gpu_pkg_op_args_t
														// removed localparam type VX_gpu_pkg_operands_t
														localparam OUT_DATAW = 473;
														// Trace: src/VX_opc_unit.sv:24:5
														wire [2:0] src_valid;
														// Trace: src/VX_opc_unit.sv:25:5
														wire [2:0] req_valid_in;
														wire [2:0] req_ready_in;
														// Trace: src/VX_opc_unit.sv:26:5
														wire [8:0] req_addr_in;
														// Trace: src/VX_opc_unit.sv:27:5
														wire [5:0] req_bank_idx;
														// Trace: src/VX_opc_unit.sv:28:5
														wire [3:0] gpr_rd_valid;
														wire [3:0] gpr_rd_ready;
														// Trace: src/VX_opc_unit.sv:29:5
														wire [3:0] gpr_rd_valid_st1;
														wire [3:0] gpr_rd_valid_st2;
														// Trace: src/VX_opc_unit.sv:30:5
														wire [11:0] gpr_rd_reg;
														wire [11:0] gpr_rd_reg_st1;
														// Trace: src/VX_opc_unit.sv:31:5
														wire [511:0] gpr_rd_data_st2;
														// Trace: src/VX_opc_unit.sv:32:5
														wire [7:0] gpr_rd_opd;
														wire [7:0] gpr_rd_opd_st1;
														wire [7:0] gpr_rd_opd_st2;
														// Trace: src/VX_opc_unit.sv:33:5
														wire [3:0] simd_out;
														// Trace: src/VX_opc_unit.sv:34:5
														wire [0:0] simd_pid;
														// Trace: src/VX_opc_unit.sv:35:5
														wire simd_sop;
														wire simd_eop;
														// Trace: src/VX_opc_unit.sv:36:5
														wire pipe_ready_in;
														// Trace: src/VX_opc_unit.sv:37:5
														wire pipe_valid_st1;
														wire pipe_ready_st1;
														// Trace: src/VX_opc_unit.sv:38:5
														wire pipe_valid_st2;
														wire pipe_ready_st2;
														// Trace: src/VX_opc_unit.sv:39:5
														wire [88:0] pipe_mdata;
														wire [88:0] pipe_mdata_st1;
														wire [88:0] pipe_mdata_st2;
														// Trace: src/VX_opc_unit.sv:40:5
														reg [383:0] opd_buffer_st2;
														reg [383:0] opd_buffer_n_st2;
														// Trace: src/VX_opc_unit.sv:41:5
														reg [2:0] opd_fetched_st1;
														// Trace: src/VX_opc_unit.sv:42:5
														reg has_collision;
														// Trace: src/VX_opc_unit.sv:43:5
														wire has_collision_st1;
														// Trace: src/VX_opc_unit.sv:44:5
														wire [14:0] src_regs;
														// Trace: src/VX_opc_unit.sv:45:5
														localparam VX_gpu_pkg_REG_TYPE_BITS = 1;
														localparam VX_gpu_pkg_RV_REGS_BITS = 5;
														// removed localparam type VX_gpu_pkg_reg_idx_t
														function automatic [4:0] VX_gpu_pkg_to_reg_number;
															// Trace: src/VX_gpu_pkg.sv:592:64
															input reg [5:0] reg_idx;
															// Trace: src/VX_gpu_pkg.sv:593:9
															VX_gpu_pkg_to_reg_number = reg_idx[4-:5];
														endfunction
														assign src_regs = {VX_gpu_pkg_to_reg_number(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[5-:6]), VX_gpu_pkg_to_reg_number(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[11-:6]), VX_gpu_pkg_to_reg_number(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[17-:6])};
														// Trace: src/VX_opc_unit.sv:48:5
														genvar _gv_i_1;
														for (_gv_i_1 = 0; _gv_i_1 < VX_gpu_pkg_NUM_SRC_OPDS; _gv_i_1 = _gv_i_1 + 1) begin : g_gpr_rd_reg
															localparam i = _gv_i_1;
															// Trace: src/VX_opc_unit.sv:49:9
															assign req_addr_in[i * 3+:3] = src_regs[(i * 5) + 4-:REG_REM_BITS];
														end
														// Trace: src/VX_opc_unit.sv:51:5
														genvar _gv_i_2;
														for (_gv_i_2 = 0; _gv_i_2 < VX_gpu_pkg_NUM_SRC_OPDS; _gv_i_2 = _gv_i_2 + 1) begin : g_req_bank_idx
															localparam i = _gv_i_2;
															if (1) begin : g_bn
																// Trace: src/VX_opc_unit.sv:53:13
																assign req_bank_idx[i * 2+:2] = src_regs[(i * 5) + 1-:2];
															end
														end
														// Trace: src/VX_opc_unit.sv:58:5
														genvar _gv_i_3;
														for (_gv_i_3 = 0; _gv_i_3 < VX_gpu_pkg_NUM_SRC_OPDS; _gv_i_3 = _gv_i_3 + 1) begin : g_src_valid
															localparam i = _gv_i_3;
															// Trace: src/VX_opc_unit.sv:59:9
															assign src_valid[i] = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[24 + i] && (src_regs[i * 5+:5] != 0)) && ~opd_fetched_st1[i];
														end
														// Trace: src/VX_opc_unit.sv:61:5
														assign req_valid_in = {VX_gpu_pkg_NUM_SRC_OPDS {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.valid}} & src_valid;
														// Trace: src/VX_opc_unit.sv:62:5
														VX_stream_xbar #(
															.NUM_INPUTS(VX_gpu_pkg_NUM_SRC_OPDS),
															.NUM_OUTPUTS(NUM_BANKS),
															.DATAW(REG_REM_BITS),
															.ARBITER("P"),
															.OUT_BUF(0)
														) req_xbar(
															.clk(clk),
															.reset(reset),
															.collisions(),
															.valid_in(req_valid_in),
															.data_in(req_addr_in),
															.sel_in(req_bank_idx),
															.ready_in(req_ready_in),
															.valid_out(gpr_rd_valid),
															.data_out(gpr_rd_reg),
															.sel_out(gpr_rd_opd),
															.ready_out(gpr_rd_ready)
														);
														// Trace: src/VX_opc_unit.sv:81:5
														assign gpr_rd_ready = {NUM_BANKS {pipe_ready_in}};
														// Trace: src/VX_opc_unit.sv:82:5
														always @(*) begin
															// Trace: src/VX_opc_unit.sv:83:9
															has_collision = 0;
															// Trace: src/VX_opc_unit.sv:84:9
															begin : sv2v_autoblock_5
																// Trace: src/VX_opc_unit.sv:84:14
																integer i;
																// Trace: src/VX_opc_unit.sv:84:14
																for (i = 0; i < VX_gpu_pkg_NUM_SRC_OPDS; i = i + 1)
																	begin
																		// Trace: src/VX_opc_unit.sv:85:13
																		begin : sv2v_autoblock_6
																			// Trace: src/VX_opc_unit.sv:85:18
																			integer j;
																			// Trace: src/VX_opc_unit.sv:85:18
																			for (j = 1; j < (VX_gpu_pkg_NUM_SRC_OPDS - i); j = j + 1)
																				begin
																					// Trace: src/VX_opc_unit.sv:86:17
																					has_collision = has_collision | ((src_valid[i] && src_valid[j + i]) && (req_bank_idx[i * 2+:2] == req_bank_idx[(j + i) * 2+:2]));
																				end
																		end
																	end
															end
														end
														// Trace: src/VX_opc_unit.sv:92:5
														wire opd_last_fetch = pipe_ready_in && ~has_collision;
														// Trace: src/VX_opc_unit.sv:93:5
														VX_nz_iterator #(
															.DATAW(4),
															.N(VX_gpu_pkg_SIMD_COUNT)
														) simd_iter(
															.clk(clk),
															.reset(reset),
															.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.valid),
															.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[104-:4]),
															.next(opd_last_fetch),
															.valid_out(),
															.data_out(simd_out),
															.pid(simd_pid),
															.sop(simd_sop),
															.eop(simd_eop)
														);
														// Trace: src/VX_opc_unit.sv:108:5
														assign pipe_mdata = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[107], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[106-:2], simd_pid, simd_out, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[100-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[27], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[70-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[68-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[64-:37], VX_gpu_pkg_to_reg_number(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.data[23-:6]), simd_sop, simd_eop};
														// Trace: src/VX_opc_unit.sv:122:5
														assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.ready = opd_last_fetch && simd_eop;
														// Trace: src/VX_opc_unit.sv:123:5
														wire pipe_fire_st1 = pipe_valid_st1 && pipe_ready_st1;
														// Trace: src/VX_opc_unit.sv:124:5
														wire pipe_fire_st2 = pipe_valid_st2 && pipe_ready_st2;
														// Trace: src/VX_opc_unit.sv:125:5
														VX_pipe_buffer #(
															.DATAW(114),
															.RESETW(1)
														) pipe_reg1(
															.clk(clk),
															.reset(reset),
															.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_scoreboard_if.valid),
															.ready_in(pipe_ready_in),
															.data_in({gpr_rd_valid, pipe_mdata, has_collision, gpr_rd_reg, gpr_rd_opd}),
															.data_out({gpr_rd_valid_st1, pipe_mdata_st1, has_collision_st1, gpr_rd_reg_st1, gpr_rd_opd_st1}),
															.valid_out(pipe_valid_st1),
															.ready_out(pipe_ready_st1)
														);
														// Trace: src/VX_opc_unit.sv:138:5
														wire [2:0] req_fire_in = req_valid_in & req_ready_in;
														// Trace: src/VX_opc_unit.sv:139:5
														always @(posedge clk)
															// Trace: src/VX_opc_unit.sv:140:9
															if (reset || opd_last_fetch)
																// Trace: src/VX_opc_unit.sv:141:13
																opd_fetched_st1 <= 1'sb0;
															else
																// Trace: src/VX_opc_unit.sv:143:13
																opd_fetched_st1 <= opd_fetched_st1 | req_fire_in;
														// Trace: src/VX_opc_unit.sv:146:5
														wire pipe_valid2_st1 = pipe_valid_st1 && ~has_collision_st1;
														// Trace: src/VX_opc_unit.sv:147:5
														VX_pipe_buffer #(
															.DATAW(101),
															.RESETW(1)
														) pipe_reg2(
															.clk(clk),
															.reset(reset),
															.valid_in(pipe_valid2_st1),
															.ready_in(pipe_ready_st1),
															.data_in({gpr_rd_valid_st1, gpr_rd_opd_st1, pipe_mdata_st1}),
															.data_out({gpr_rd_valid_st2, gpr_rd_opd_st2, pipe_mdata_st2}),
															.valid_out(pipe_valid_st2),
															.ready_out(pipe_ready_st2)
														);
														// Trace: src/VX_opc_unit.sv:160:5
														always @(*) begin
															// Trace: src/VX_opc_unit.sv:161:9
															opd_buffer_n_st2 = opd_buffer_st2;
															// Trace: src/VX_opc_unit.sv:162:9
															begin : sv2v_autoblock_7
																// Trace: src/VX_opc_unit.sv:162:14
																integer b;
																// Trace: src/VX_opc_unit.sv:162:14
																for (b = 0; b < NUM_BANKS; b = b + 1)
																	begin
																		// Trace: src/VX_opc_unit.sv:163:13
																		if (gpr_rd_valid_st2[b])
																			// Trace: src/VX_opc_unit.sv:164:17
																			opd_buffer_n_st2[gpr_rd_opd_st2[b * 2+:2] * 128+:128] = gpr_rd_data_st2[32 * (b * 4)+:128];
																	end
															end
														end
														// Trace: src/VX_opc_unit.sv:168:5
														always @(posedge clk)
															// Trace: src/VX_opc_unit.sv:169:9
															if (reset || pipe_fire_st2)
																// Trace: src/VX_opc_unit.sv:170:13
																opd_buffer_st2 <= 1'sb0;
															else
																// Trace: src/VX_opc_unit.sv:172:13
																opd_buffer_st2 <= opd_buffer_n_st2;
														// Trace: src/VX_opc_unit.sv:175:5
														wire [4:0] gpr_wr_addr;
														// Trace: src/VX_opc_unit.sv:176:5
														if (1) begin : g_gpr_wr_addr
															if (1) begin : genblk1
																// Trace: src/VX_opc_unit.sv:195:9
																assign gpr_wr_addr = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_writeback_if.data[171-:PER_OPC_NW_BITS], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_writeback_if.data[134-:REG_REM_BITS]};
															end
														end
														// Trace: src/VX_opc_unit.sv:199:5
														wire [1:0] gpr_wr_bank_idx;
														// Trace: src/VX_opc_unit.sv:200:5
														if (1) begin : g_gpr_wr_bank_idx_bn
															// Trace: src/VX_opc_unit.sv:201:9
															assign gpr_wr_bank_idx = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_writeback_if.data[131:130];
														end
														// Trace: src/VX_opc_unit.sv:205:5
														wire [15:0] gpr_wr_byteen;
														// Trace: src/VX_opc_unit.sv:206:5
														genvar _gv_i_4;
														localparam VX_gpu_pkg_XLENB = 4;
														for (_gv_i_4 = 0; _gv_i_4 < 4; _gv_i_4 = _gv_i_4 + 1) begin : g_gpr_wr_byteen
															localparam i = _gv_i_4;
															// Trace: src/VX_opc_unit.sv:207:9
															assign gpr_wr_byteen[i * VX_gpu_pkg_XLENB+:VX_gpu_pkg_XLENB] = {VX_gpu_pkg_XLENB {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_writeback_if.data[165 + i]}};
														end
														// Trace: src/VX_opc_unit.sv:209:5
														genvar _gv_b_1;
														for (_gv_b_1 = 0; _gv_b_1 < NUM_BANKS; _gv_b_1 = _gv_b_1 + 1) begin : g_gpr_rams
															localparam b = _gv_b_1;
															// Trace: src/VX_opc_unit.sv:210:9
															wire gpr_wr_enabled;
															if (1) begin : g_gpr_wr_enabled_bn
																// Trace: src/VX_opc_unit.sv:212:13
																assign gpr_wr_enabled = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_writeback_if.valid && (gpr_wr_bank_idx == sv2v_cast_2_signed(b));
															end
															// Trace: src/VX_opc_unit.sv:216:9
															wire [4:0] gpr_rd_addr;
															if (1) begin : g_gpr_rd_addr
																if (1) begin : genblk1
																	// Trace: src/VX_opc_unit.sv:236:9
																	assign gpr_rd_addr = {pipe_mdata_st1[87-:PER_OPC_NW_BITS], gpr_rd_reg_st1[b * 3+:3]};
																end
															end
															// Trace: src/VX_opc_unit.sv:240:9
															VX_dp_ram #(
																.DATAW(BANK_DATA_WIDTH),
																.SIZE(BANK_SIZE),
																.WRENW(BANK_DATA_SIZE),
																.OUT_REG(1),
																.RDW_MODE("R")
															) gpr_ram(
																.clk(clk),
																.reset(reset),
																.read(pipe_fire_st1),
																.wren(gpr_wr_byteen),
																.write(gpr_wr_enabled),
																.waddr(gpr_wr_addr),
																.wdata(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.g_collectors[_gv_i_206].opc_writeback_if.data[129-:128]),
																.raddr(gpr_rd_addr),
																.rdata(gpr_rd_data_st2[32 * (b * 4)+:128])
															);
														end
														// Trace: src/VX_opc_unit.sv:258:5
														VX_elastic_buffer #(
															.DATAW(OUT_DATAW),
															.SIZE(2),
															.OUT_REG(1)
														) out_buf(
															.clk(clk),
															.reset(reset),
															.valid_in(pipe_valid_st2),
															.ready_in(pipe_ready_st2),
															.data_in({pipe_mdata_st2[88:2], opd_buffer_n_st2, pipe_mdata_st2[1:0]}),
															.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[472], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[471-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[469], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[468-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[464-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[391], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[434-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[432-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[428-:37], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[390-:5], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[129-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[257-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[385-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].data[0]}),
															.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].valid),
															.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands.per_opc_operands_if[_mbase_operands_if].ready)
														);
													end
													assign opc_unit.clk = clk;
													assign opc_unit.reset = reset;
												end
												// Trace: src/VX_operands.sv:44:5
												wire [0:0] per_opc_operands_valid;
												// Trace: src/VX_operands.sv:45:5
												wire [472:0] per_opc_operands_data;
												// Trace: src/VX_operands.sv:46:5
												wire [0:0] per_opc_operands_ready;
												// Trace: src/VX_operands.sv:48:5
												genvar _gv_i_207;
												for (_gv_i_207 = 0; _gv_i_207 < 1; _gv_i_207 = _gv_i_207 + 1) begin : genblk3
													localparam i = _gv_i_207;
													// Trace: src/VX_operands.sv:49:9
													assign per_opc_operands_valid[i] = per_opc_operands_if[i].valid;
													// Trace: src/VX_operands.sv:50:9
													assign per_opc_operands_data[i * 473+:473] = per_opc_operands_if[i].data;
													// Trace: src/VX_operands.sv:51:9
													assign per_opc_operands_if[i].ready = per_opc_operands_ready[i];
												end
												// Trace: src/VX_operands.sv:54:5
												VX_stream_arb #(
													.NUM_INPUTS(1),
													.NUM_OUTPUTS(1),
													.DATAW(OUT_DATAW),
													.ARBITER("P"),
													.STICKY(OUT_ARB_STICKY),
													.OUT_BUF(0)
												) output_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(per_opc_operands_valid),
													.data_in(per_opc_operands_data),
													.ready_in(per_opc_operands_ready),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.valid),
													.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.ready),
													.sel_out()
												);
											end
											assign operands.clk = clk;
											assign operands.reset = reset;
											// Trace: src/VX_issue_slice.sv:44:5
											// expanded module instance: dispatch
											localparam _bbase_1A128_dispatch_if = 0;
											localparam _param_1A128_INSTANCE_ID = "";
											localparam _param_1A128_ISSUE_ID = ISSUE_ID;
											if (1) begin : dispatch
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_dispatch.sv:2:15
												localparam INSTANCE_ID = _param_1A128_INSTANCE_ID;
												// Trace: src/VX_dispatch.sv:3:15
												localparam ISSUE_ID = _param_1A128_ISSUE_ID;
												// Trace: src/VX_dispatch.sv:5:5
												wire clk;
												// Trace: src/VX_dispatch.sv:6:5
												wire reset;
												// Trace: src/VX_dispatch.sv:7:5
												// removed modport instance operands_if
												// Trace: src/VX_dispatch.sv:8:5
												localparam VX_gpu_pkg_EX_SFU = 2;
												localparam VX_gpu_pkg_EX_FPU = 2;
												localparam VX_gpu_pkg_EX_TCU = 2;
												localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
												localparam _mbase_dispatch_if = 0;
												// Trace: src/VX_dispatch.sv:10:5
												localparam VX_gpu_pkg_INST_ALU_BITS = 4;
												localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
												localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
												localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_RV_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
												localparam VX_gpu_pkg_PC_BITS = 30;
												localparam VX_gpu_pkg_SIMD_COUNT = 1;
												localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
												localparam VX_gpu_pkg_SIMD_IDX_W = 1;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
												// removed localparam type VX_gpu_pkg_alu_args_t
												localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
												// removed localparam type VX_gpu_pkg_csr_args_t
												localparam VX_gpu_pkg_INST_FMT_BITS = 2;
												localparam VX_gpu_pkg_INST_FRM_BITS = 3;
												// removed localparam type VX_gpu_pkg_fpu_args_t
												localparam VX_gpu_pkg_OFFSET_BITS = 12;
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												// removed localparam type VX_gpu_pkg_dispatch_t
												localparam OUT_DATAW = 471;
												// Trace: src/VX_dispatch.sv:11:5
												wire [2:0] operands_ready_in;
												// Trace: src/VX_dispatch.sv:12:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.ready = operands_ready_in[Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[434-:2]];
												// Trace: src/VX_dispatch.sv:13:5
												genvar _gv_i_91;
												localparam VX_gpu_pkg_EX_BITS = 2;
												for (_gv_i_91 = 0; _gv_i_91 < VX_gpu_pkg_NUM_EX_UNITS; _gv_i_91 = _gv_i_91 + 1) begin : g_buffers
													localparam i = _gv_i_91;
													// Trace: src/VX_dispatch.sv:14:9
													VX_elastic_buffer #(
														.DATAW(OUT_DATAW),
														.SIZE(2),
														.OUT_REG(1)
													) buffer(
														.clk(clk),
														.reset(reset),
														.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.valid && (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[434-:2] == sv2v_cast_2_signed(i))),
														.ready_in(operands_ready_in[i]),
														.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[472], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[471-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[469], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[468-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[464-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[432-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[428-:37], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[391], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[390-:5], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[385-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[257-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[129-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].issue_slice.operands_if.data[0]}),
														.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_dispatch_if[i + _mbase_dispatch_if].data),
														.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_dispatch_if[i + _mbase_dispatch_if].valid),
														.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue.g_slices[_gv_issue_id_1].per_issue_dispatch_if[i + _mbase_dispatch_if].ready)
													);
												end
											end
											assign dispatch.clk = clk;
											assign dispatch.reset = reset;
											// Trace: src/VX_issue_slice.sv:53:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue_sched_if[_mbase_issue_sched_if].valid = (operands_if.valid && operands_if.ready) && operands_if.data[1];
											// Trace: src/VX_issue_slice.sv:54:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.issue_sched_if[_mbase_issue_sched_if].wis = operands_if.data[471-:2];
										end
										assign issue_slice.clk = clk;
										assign issue_slice.reset = reset;
										genvar _gv_ex_id_1;
										for (_gv_ex_id_1 = 0; _gv_ex_id_1 < VX_gpu_pkg_NUM_EX_UNITS; _gv_ex_id_1 = _gv_ex_id_1 + 1) begin : g_dispatch_if
											localparam ex_id = _gv_ex_id_1;
											// Trace: src/VX_issue.sv:33:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[((ex_id * 1) + issue_id) + _mbase_dispatch_if].valid = per_issue_dispatch_if[ex_id].valid;
											// Trace: src/VX_issue.sv:34:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[((ex_id * 1) + issue_id) + _mbase_dispatch_if].data = per_issue_dispatch_if[ex_id].data;
											// Trace: src/VX_issue.sv:35:5
											assign per_issue_dispatch_if[ex_id].ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[((ex_id * 1) + issue_id) + _mbase_dispatch_if].ready;
										end
									end
								end
								assign issue.clk = clk;
								assign issue.reset = reset;
								// Trace: src/VX_core.sv:82:5
								// expanded module instance: execute
								localparam _bbase_B78CA_lsu_mem_if = 0;
								localparam _bbase_B78CA_dispatch_if = 0;
								localparam _bbase_B78CA_commit_if = 0;
								localparam _bbase_B78CA_branch_ctl_if = 0;
								localparam _param_B78CA_INSTANCE_ID = "";
								localparam _param_B78CA_CORE_ID = CORE_ID;
								if (1) begin : execute
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_execute.sv:2:15
									localparam INSTANCE_ID = _param_B78CA_INSTANCE_ID;
									// Trace: src/VX_execute.sv:3:15
									localparam CORE_ID = _param_B78CA_CORE_ID;
									// Trace: src/VX_execute.sv:5:5
									wire clk;
									// Trace: src/VX_execute.sv:6:5
									wire reset;
									// Trace: src/VX_execute.sv:7:5
									// removed localparam type VX_gpu_pkg_base_dcrs_t
									wire [71:0] base_dcrs;
									// Trace: src/VX_execute.sv:8:5
									localparam _mbase_lsu_mem_if = 0;
									// Trace: src/VX_execute.sv:9:5
									localparam VX_gpu_pkg_EX_SFU = 2;
									localparam VX_gpu_pkg_EX_FPU = 2;
									localparam VX_gpu_pkg_EX_TCU = 2;
									localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
									localparam _mbase_dispatch_if = 0;
									// Trace: src/VX_execute.sv:10:5
									localparam _mbase_commit_if = 0;
									// Trace: src/VX_execute.sv:11:5
									// removed modport instance sched_csr_if
									// Trace: src/VX_execute.sv:12:5
									localparam _mbase_branch_ctl_if = 0;
									// Trace: src/VX_execute.sv:13:5
									// removed modport instance warp_ctl_if
									// Trace: src/VX_execute.sv:14:5
									// removed modport instance commit_csr_if
									// Trace: src/VX_execute.sv:16:5
									localparam VX_gpu_pkg_EX_ALU = 0;
									// expanded module instance: alu_unit
									localparam _bbase_4B10A_dispatch_if = 0;
									localparam _bbase_4B10A_commit_if = 0;
									localparam _bbase_4B10A_branch_ctl_if = 0;
									localparam _param_4B10A_INSTANCE_ID = "";
									if (1) begin : alu_unit
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_alu_unit.sv:2:15
										localparam INSTANCE_ID = _param_4B10A_INSTANCE_ID;
										// Trace: src/VX_alu_unit.sv:4:5
										wire clk;
										// Trace: src/VX_alu_unit.sv:5:5
										wire reset;
										// Trace: src/VX_alu_unit.sv:6:5
										localparam _mbase_dispatch_if = 0;
										// Trace: src/VX_alu_unit.sv:7:5
										localparam _mbase_commit_if = 0;
										// Trace: src/VX_alu_unit.sv:8:5
										localparam _mbase_branch_ctl_if = 0;
										// Trace: src/VX_alu_unit.sv:10:5
										localparam BLOCK_SIZE = 1;
										// Trace: src/VX_alu_unit.sv:11:5
										localparam NUM_LANES = 4;
										// Trace: src/VX_alu_unit.sv:12:5
										localparam PARTIAL_BW = 1'd0;
										// Trace: src/VX_alu_unit.sv:13:5
										localparam PE_COUNT = 2;
										// Trace: src/VX_alu_unit.sv:14:5
										localparam PE_SEL_BITS = 1;
										// Trace: src/VX_alu_unit.sv:15:5
										localparam PE_IDX_INT = 0;
										// Trace: src/VX_alu_unit.sv:16:5
										localparam PE_IDX_MDV = 1;
										// Trace: src/VX_alu_unit.sv:17:5
										// expanded interface instance: per_block_execute_if
										localparam _param_E2592_NUM_LANES = NUM_LANES;
										genvar _arr_E2592;
										for (_arr_E2592 = 0; _arr_E2592 <= 0; _arr_E2592 = _arr_E2592 + 1) begin : per_block_execute_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_execute_if.sv:2:15
											localparam NUM_LANES = _param_E2592_NUM_LANES;
											// Trace: src/VX_execute_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_execute_if.sv:5:5
											localparam VX_gpu_pkg_INST_ALU_BITS = 4;
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
											// removed localparam type VX_gpu_pkg_alu_args_t
											localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
											// removed localparam type VX_gpu_pkg_csr_args_t
											localparam VX_gpu_pkg_INST_FMT_BITS = 2;
											localparam VX_gpu_pkg_INST_FRM_BITS = 3;
											// removed localparam type VX_gpu_pkg_fpu_args_t
											localparam VX_gpu_pkg_OFFSET_BITS = 12;
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											// removed localparam type data_t
											// Trace: src/VX_execute_if.sv:21:5
											wire valid;
											// Trace: src/VX_execute_if.sv:22:5
											wire [470:0] data;
											// Trace: src/VX_execute_if.sv:23:5
											wire ready;
											// Trace: src/VX_execute_if.sv:24:5
											// Trace: src/VX_execute_if.sv:29:5
										end
										// Trace: src/VX_alu_unit.sv:20:5
										// expanded interface instance: per_block_result_if
										localparam _param_911F6_NUM_LANES = NUM_LANES;
										genvar _arr_911F6;
										for (_arr_911F6 = 0; _arr_911F6 <= 0; _arr_911F6 = _arr_911F6 + 1) begin : per_block_result_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_result_if.sv:2:15
											localparam NUM_LANES = _param_911F6_NUM_LANES;
											// Trace: src/VX_result_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_result_if.sv:5:5
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											// removed localparam type data_t
											// Trace: src/VX_result_if.sv:17:5
											wire valid;
											// Trace: src/VX_result_if.sv:18:5
											wire [173:0] data;
											// Trace: src/VX_result_if.sv:19:5
											wire ready;
											// Trace: src/VX_result_if.sv:20:5
											// Trace: src/VX_result_if.sv:25:5
										end
										// Trace: src/VX_alu_unit.sv:23:5
										// expanded module instance: dispatch_unit
										localparam _bbase_2E16E_dispatch_if = 0;
										localparam _bbase_2E16E_execute_if = 0;
										localparam _param_2E16E_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_2E16E_NUM_LANES = NUM_LANES;
										localparam _param_2E16E_OUT_BUF = (PARTIAL_BW ? 3 : 0);
										if (1) begin : dispatch_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_dispatch_unit.sv:2:15
											localparam BLOCK_SIZE = _param_2E16E_BLOCK_SIZE;
											// Trace: src/VX_dispatch_unit.sv:3:15
											localparam NUM_LANES = _param_2E16E_NUM_LANES;
											// Trace: src/VX_dispatch_unit.sv:4:15
											localparam OUT_BUF = _param_2E16E_OUT_BUF;
											// Trace: src/VX_dispatch_unit.sv:5:15
											localparam MAX_FANOUT = 8;
											// Trace: src/VX_dispatch_unit.sv:7:5
											wire clk;
											// Trace: src/VX_dispatch_unit.sv:8:5
											wire reset;
											// Trace: src/VX_dispatch_unit.sv:9:5
											localparam _mbase_dispatch_if = 0;
											// Trace: src/VX_dispatch_unit.sv:10:5
											localparam _mbase_execute_if = 0;
											// Trace: src/VX_dispatch_unit.sv:12:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:13:5
											localparam NUM_PACKETS = 1;
											// Trace: src/VX_dispatch_unit.sv:14:5
											localparam LPID_BITS = 0;
											// Trace: src/VX_dispatch_unit.sv:15:5
											localparam LPID_WIDTH = 1;
											// Trace: src/VX_dispatch_unit.sv:16:5
											localparam GPID_BITS = 0;
											// Trace: src/VX_dispatch_unit.sv:17:5
											localparam GPID_WIDTH = 1;
											// Trace: src/VX_dispatch_unit.sv:18:5
											localparam BATCH_COUNT = 1;
											// Trace: src/VX_dispatch_unit.sv:19:5
											localparam BATCH_COUNT_W = 1;
											// Trace: src/VX_dispatch_unit.sv:20:5
											localparam ISSUE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:21:5
											localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
											localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
											localparam VX_gpu_pkg_INST_OP_BITS = 4;
											localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
											localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
											localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_SIMD_COUNT = 1;
											localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
											localparam VX_gpu_pkg_SIMD_IDX_W = 1;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam IN_DATAW = 471;
											// Trace: src/VX_dispatch_unit.sv:22:5
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam OUT_DATAW = 471;
											// Trace: src/VX_dispatch_unit.sv:23:5
											localparam FANOUT_ENABLE = 1'd0;
											// Trace: src/VX_dispatch_unit.sv:24:5
											localparam DATA_TMASK_OFF = 463;
											// Trace: src/VX_dispatch_unit.sv:25:5
											localparam DATA_REGS_OFF = 2;
											// Trace: src/VX_dispatch_unit.sv:26:5
											// removed localparam type packet_t
											// Trace: src/VX_dispatch_unit.sv:30:5
											wire [0:0] dispatch_valid;
											// Trace: src/VX_dispatch_unit.sv:31:5
											wire [470:0] dispatch_data;
											// Trace: src/VX_dispatch_unit.sv:32:5
											wire [0:0] dispatch_ready;
											// Trace: src/VX_dispatch_unit.sv:33:5
											genvar _gv_i_35;
											for (_gv_i_35 = 0; _gv_i_35 < 1; _gv_i_35 = _gv_i_35 + 1) begin : g_dispatch_data
												localparam i = _gv_i_35;
												// Trace: src/VX_dispatch_unit.sv:34:9
												assign dispatch_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].valid;
												// Trace: src/VX_dispatch_unit.sv:35:9
												assign dispatch_data[i * 471+:471] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].data;
												// Trace: src/VX_dispatch_unit.sv:36:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].ready = dispatch_ready[i];
											end
											// Trace: src/VX_dispatch_unit.sv:38:5
											wire [0:0] block_ready;
											// Trace: src/VX_dispatch_unit.sv:39:5
											wire [3:0] block_tmask;
											// Trace: src/VX_dispatch_unit.sv:40:5
											wire [383:0] block_rsdata;
											// Trace: src/VX_dispatch_unit.sv:41:5
											wire [0:0] block_pid;
											// Trace: src/VX_dispatch_unit.sv:42:5
											wire [0:0] block_sop;
											// Trace: src/VX_dispatch_unit.sv:43:5
											wire [0:0] block_eop;
											// Trace: src/VX_dispatch_unit.sv:44:5
											wire [0:0] block_done;
											// Trace: src/VX_dispatch_unit.sv:45:5
											wire batch_done = &block_done;
											// Trace: src/VX_dispatch_unit.sv:46:5
											wire [0:0] batch_idx;
											// Trace: src/VX_dispatch_unit.sv:47:5
											if (1) begin : g_batch_idx_0
												// Trace: src/VX_dispatch_unit.sv:73:9
												assign batch_idx = 0;
											end
											// Trace: src/VX_dispatch_unit.sv:75:5
											wire [0:0] issue_indices;
											// Trace: src/VX_dispatch_unit.sv:76:5
											genvar _gv_block_idx_2;
											for (_gv_block_idx_2 = 0; _gv_block_idx_2 < BLOCK_SIZE; _gv_block_idx_2 = _gv_block_idx_2 + 1) begin : g_issue_indices
												localparam block_idx = _gv_block_idx_2;
												// Trace: src/VX_dispatch_unit.sv:77:9
												assign issue_indices[block_idx+:1] = sv2v_cast_1(batch_idx * BLOCK_SIZE) + sv2v_cast_1_signed(block_idx);
											end
											// Trace: src/VX_dispatch_unit.sv:79:5
											genvar _gv_block_idx_3;
											localparam VX_gpu_pkg_ISSUE_ISW_BITS = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											function automatic [1:0] VX_gpu_pkg_wis_to_wid;
												// Trace: src/VX_gpu_pkg.sv:264:9
												input reg [1:0] wis;
												// Trace: src/VX_gpu_pkg.sv:265:9
												input reg [0:0] isw;
												// Trace: src/VX_gpu_pkg.sv:267:9
												begin
													// Trace: src/VX_gpu_pkg.sv:270:13
													VX_gpu_pkg_wis_to_wid = wis;
												end
											endfunction
											for (_gv_block_idx_3 = 0; _gv_block_idx_3 < BLOCK_SIZE; _gv_block_idx_3 = _gv_block_idx_3 + 1) begin : g_blocks
												localparam block_idx = _gv_block_idx_3;
												// Trace: src/VX_dispatch_unit.sv:80:9
												wire [0:0] issue_idx = issue_indices[block_idx+:1];
												// Trace: src/VX_dispatch_unit.sv:81:9
												wire [1:0] dispatch_wis = dispatch_data[(issue_idx * 471) + 468+:VX_gpu_pkg_ISSUE_WIS_W];
												// Trace: src/VX_dispatch_unit.sv:82:9
												wire [0:0] dispatch_sid = dispatch_data[(issue_idx * 471) + 467+:VX_gpu_pkg_SIMD_IDX_W];
												// Trace: src/VX_dispatch_unit.sv:83:9
												wire dispatch_sop = dispatch_data[(issue_idx * 471) + 1];
												// Trace: src/VX_dispatch_unit.sv:84:9
												wire dispatch_eop = dispatch_data[issue_idx * 471];
												// Trace: src/VX_dispatch_unit.sv:85:9
												wire [3:0] dispatch_tmask;
												// Trace: src/VX_dispatch_unit.sv:86:9
												wire [383:0] dispatch_rsdata;
												// Trace: src/VX_dispatch_unit.sv:87:9
												assign dispatch_tmask = dispatch_data[(issue_idx * 471) + DATA_TMASK_OFF+:4];
												// Trace: src/VX_dispatch_unit.sv:88:9
												assign dispatch_rsdata[0+:128] = dispatch_data[(issue_idx * 471) + 258+:128];
												// Trace: src/VX_dispatch_unit.sv:89:9
												assign dispatch_rsdata[128+:128] = dispatch_data[(issue_idx * 471) + 130+:128];
												// Trace: src/VX_dispatch_unit.sv:90:9
												assign dispatch_rsdata[256+:128] = dispatch_data[(issue_idx * 471) + 2+:128];
												// Trace: src/VX_dispatch_unit.sv:91:9
												wire valid_p;
												wire ready_p;
												if (1) begin : g_full_simd
													// Trace: src/VX_dispatch_unit.sv:132:13
													assign valid_p = dispatch_valid[issue_idx];
													// Trace: src/VX_dispatch_unit.sv:133:13
													assign block_tmask[block_idx * 4+:4] = dispatch_tmask;
													// Trace: src/VX_dispatch_unit.sv:134:13
													assign block_rsdata[32 * (4 * (block_idx * 3))+:384] = dispatch_rsdata;
													// Trace: src/VX_dispatch_unit.sv:135:13
													assign block_pid[block_idx+:1] = 0;
													// Trace: src/VX_dispatch_unit.sv:136:13
													assign block_sop[block_idx] = 1;
													// Trace: src/VX_dispatch_unit.sv:137:13
													assign block_eop[block_idx] = 1;
													// Trace: src/VX_dispatch_unit.sv:138:13
													assign block_ready[block_idx] = ready_p;
													// Trace: src/VX_dispatch_unit.sv:139:13
													assign block_done[block_idx] = ready_p || ~valid_p;
												end
												// Trace: src/VX_dispatch_unit.sv:141:9
												wire [0:0] isw;
												if (1) begin : g_isw
													// Trace: src/VX_dispatch_unit.sv:149:13
													assign isw = block_idx;
												end
												// Trace: src/VX_dispatch_unit.sv:151:9
												wire [1:0] block_wid = VX_gpu_pkg_wis_to_wid(dispatch_wis, isw);
												// Trace: src/VX_dispatch_unit.sv:152:9
												wire [0:0] warp_pid = block_pid[block_idx+:1] + sv2v_cast_1(dispatch_sid * NUM_PACKETS);
												// Trace: src/VX_dispatch_unit.sv:153:9
												wire warp_sop = block_sop[block_idx] && dispatch_sop;
												// Trace: src/VX_dispatch_unit.sv:154:9
												wire warp_eop = block_eop[block_idx] && dispatch_eop;
												// Trace: src/VX_dispatch_unit.sv:155:9
												VX_elastic_buffer #(
													.DATAW(OUT_DATAW),
													.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
													.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
												) buf_out(
													.clk(clk),
													.reset(reset),
													.valid_in(valid_p),
													.ready_in(ready_p),
													.data_in({dispatch_data[(issue_idx * 471) + 470-:VX_gpu_pkg_UUID_WIDTH], block_wid, block_tmask[block_idx * 4+:4], dispatch_data[(issue_idx * 471) + 462-:77], block_rsdata[32 * ((block_idx * 3) * 4)+:128], block_rsdata[32 * (((block_idx * 3) + 1) * 4)+:128], block_rsdata[32 * (((block_idx * 3) + 2) * 4)+:128], warp_pid, warp_sop, warp_eop}),
													.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_execute_if[block_idx + _mbase_execute_if].data),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_execute_if[block_idx + _mbase_execute_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_execute_if[block_idx + _mbase_execute_if].ready)
												);
											end
											// Trace: src/VX_dispatch_unit.sv:180:5
											reg [0:0] ready_in;
											// Trace: src/VX_dispatch_unit.sv:181:5
											always @(*) begin
												// Trace: src/VX_dispatch_unit.sv:182:9
												ready_in = 0;
												// Trace: src/VX_dispatch_unit.sv:183:9
												begin : sv2v_autoblock_8
													// Trace: src/VX_dispatch_unit.sv:183:14
													integer block_idx;
													// Trace: src/VX_dispatch_unit.sv:183:14
													for (block_idx = 0; block_idx < BLOCK_SIZE; block_idx = block_idx + 1)
														begin
															// Trace: src/VX_dispatch_unit.sv:184:13
															ready_in[issue_indices[block_idx+:1]] = block_ready[block_idx] && block_eop[block_idx];
														end
												end
											end
											// Trace: src/VX_dispatch_unit.sv:187:5
											assign dispatch_ready = ready_in;
										end
										assign dispatch_unit.clk = clk;
										assign dispatch_unit.reset = reset;
										// Trace: src/VX_alu_unit.sv:33:5
										genvar _gv_block_idx_1;
										localparam VX_gpu_pkg_ALU_TYPE_MULDIV = 2;
										for (_gv_block_idx_1 = 0; _gv_block_idx_1 < BLOCK_SIZE; _gv_block_idx_1 = _gv_block_idx_1 + 1) begin : g_blocks
											localparam block_idx = _gv_block_idx_1;
											// Trace: src/VX_alu_unit.sv:34:9
											// expanded interface instance: pe_execute_if
											localparam _param_C9035_NUM_LANES = NUM_LANES;
											genvar _arr_C9035;
											for (_arr_C9035 = 0; _arr_C9035 <= 1; _arr_C9035 = _arr_C9035 + 1) begin : pe_execute_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_execute_if.sv:2:15
												localparam NUM_LANES = _param_C9035_NUM_LANES;
												// Trace: src/VX_execute_if.sv:3:15
												localparam PID_WIDTH = 1;
												// Trace: src/VX_execute_if.sv:5:5
												localparam VX_gpu_pkg_INST_ALU_BITS = 4;
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_RV_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
												localparam VX_gpu_pkg_NW_BITS = 2;
												localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
												localparam VX_gpu_pkg_PC_BITS = 30;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
												// removed localparam type VX_gpu_pkg_alu_args_t
												localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
												// removed localparam type VX_gpu_pkg_csr_args_t
												localparam VX_gpu_pkg_INST_FMT_BITS = 2;
												localparam VX_gpu_pkg_INST_FRM_BITS = 3;
												// removed localparam type VX_gpu_pkg_fpu_args_t
												localparam VX_gpu_pkg_OFFSET_BITS = 12;
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												// removed localparam type data_t
												// Trace: src/VX_execute_if.sv:21:5
												wire valid;
												// Trace: src/VX_execute_if.sv:22:5
												wire [470:0] data;
												// Trace: src/VX_execute_if.sv:23:5
												wire ready;
												// Trace: src/VX_execute_if.sv:24:5
												// Trace: src/VX_execute_if.sv:29:5
											end
											// Trace: src/VX_alu_unit.sv:37:9
											// expanded interface instance: pe_result_if
											localparam _param_FE18D_NUM_LANES = NUM_LANES;
											genvar _arr_FE18D;
											for (_arr_FE18D = 0; _arr_FE18D <= 1; _arr_FE18D = _arr_FE18D + 1) begin : pe_result_if
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_result_if.sv:2:15
												localparam NUM_LANES = _param_FE18D_NUM_LANES;
												// Trace: src/VX_result_if.sv:3:15
												localparam PID_WIDTH = 1;
												// Trace: src/VX_result_if.sv:5:5
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_RV_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
												localparam VX_gpu_pkg_NW_BITS = 2;
												localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
												localparam VX_gpu_pkg_PC_BITS = 30;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												// removed localparam type data_t
												// Trace: src/VX_result_if.sv:17:5
												wire valid;
												// Trace: src/VX_result_if.sv:18:5
												wire [173:0] data;
												// Trace: src/VX_result_if.sv:19:5
												wire ready;
												// Trace: src/VX_result_if.sv:20:5
												// Trace: src/VX_result_if.sv:25:5
											end
											// Trace: src/VX_alu_unit.sv:40:9
											reg [0:0] pe_select;
											// Trace: src/VX_alu_unit.sv:41:9
											always @(*) begin
												// Trace: src/VX_alu_unit.sv:42:13
												pe_select = PE_IDX_INT;
												// Trace: src/VX_alu_unit.sv:43:13
												if (per_block_execute_if[block_idx].data[426-:2] == VX_gpu_pkg_ALU_TYPE_MULDIV)
													// Trace: src/VX_alu_unit.sv:44:17
													pe_select = PE_IDX_MDV;
											end
											// Trace: src/VX_alu_unit.sv:46:9
											// expanded module instance: pe_switch
											localparam _bbase_3D12E_execute_in_if = block_idx;
											localparam _bbase_3D12E_result_out_if = block_idx;
											localparam _bbase_3D12E_execute_out_if = 0;
											localparam _bbase_3D12E_result_in_if = 0;
											localparam _param_3D12E_PE_COUNT = PE_COUNT;
											localparam _param_3D12E_NUM_LANES = NUM_LANES;
											localparam _param_3D12E_ARBITER = "R";
											localparam _param_3D12E_REQ_OUT_BUF = 0;
											localparam _param_3D12E_RSP_OUT_BUF = (PARTIAL_BW ? 1 : 3);
											if (1) begin : pe_switch
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_pe_switch.sv:2:15
												localparam PE_COUNT = _param_3D12E_PE_COUNT;
												// Trace: src/VX_pe_switch.sv:3:15
												localparam NUM_LANES = _param_3D12E_NUM_LANES;
												// Trace: src/VX_pe_switch.sv:4:15
												localparam REQ_OUT_BUF = _param_3D12E_REQ_OUT_BUF;
												// Trace: src/VX_pe_switch.sv:5:15
												localparam RSP_OUT_BUF = _param_3D12E_RSP_OUT_BUF;
												// Trace: src/VX_pe_switch.sv:6:15
												localparam ARBITER = _param_3D12E_ARBITER;
												// Trace: src/VX_pe_switch.sv:7:15
												localparam PE_SEL_BITS = 1;
												// Trace: src/VX_pe_switch.sv:9:5
												wire clk;
												// Trace: src/VX_pe_switch.sv:10:5
												wire reset;
												// Trace: src/VX_pe_switch.sv:11:5
												wire [0:0] pe_sel;
												// Trace: src/VX_pe_switch.sv:12:5
												localparam _mbase_execute_in_if = _bbase_3D12E_execute_in_if;
												// Trace: src/VX_pe_switch.sv:13:5
												localparam _mbase_result_out_if = _bbase_3D12E_result_out_if;
												// Trace: src/VX_pe_switch.sv:14:5
												localparam _mbase_execute_out_if = 0;
												// Trace: src/VX_pe_switch.sv:15:5
												localparam _mbase_result_in_if = 0;
												// Trace: src/VX_pe_switch.sv:17:5
												localparam PID_BITS = 0;
												// Trace: src/VX_pe_switch.sv:18:5
												localparam PID_WIDTH = 1;
												// Trace: src/VX_pe_switch.sv:19:5
												localparam VX_gpu_pkg_INST_ALU_BITS = 4;
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_RV_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
												localparam VX_gpu_pkg_NW_BITS = 2;
												localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
												localparam VX_gpu_pkg_PC_BITS = 30;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
												// removed localparam type VX_gpu_pkg_alu_args_t
												localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
												// removed localparam type VX_gpu_pkg_csr_args_t
												localparam VX_gpu_pkg_INST_FMT_BITS = 2;
												localparam VX_gpu_pkg_INST_FRM_BITS = 3;
												// removed localparam type VX_gpu_pkg_fpu_args_t
												localparam VX_gpu_pkg_OFFSET_BITS = 12;
												// removed localparam type VX_gpu_pkg_lsu_args_t
												// removed localparam type VX_gpu_pkg_wctl_args_t
												// removed localparam type VX_gpu_pkg_op_args_t
												localparam REQ_DATAW = 471;
												// Trace: src/VX_pe_switch.sv:20:5
												localparam RSP_DATAW = 174;
												// Trace: src/VX_pe_switch.sv:21:5
												wire [1:0] pe_req_valid;
												// Trace: src/VX_pe_switch.sv:22:5
												wire [941:0] pe_req_data;
												// Trace: src/VX_pe_switch.sv:23:5
												wire [1:0] pe_req_ready;
												// Trace: src/VX_pe_switch.sv:24:5
												VX_stream_switch #(
													.DATAW(REQ_DATAW),
													.NUM_INPUTS(1),
													.NUM_OUTPUTS(PE_COUNT),
													.OUT_BUF(REQ_OUT_BUF)
												) req_switch(
													.clk(clk),
													.reset(reset),
													.sel_in(pe_sel),
													.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_execute_if[_mbase_execute_in_if].valid),
													.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_execute_if[_mbase_execute_in_if].ready),
													.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_execute_if[_mbase_execute_in_if].data),
													.data_out(pe_req_data),
													.valid_out(pe_req_valid),
													.ready_out(pe_req_ready)
												);
												// Trace: src/VX_pe_switch.sv:40:5
												genvar _gv_i_150;
												for (_gv_i_150 = 0; _gv_i_150 < PE_COUNT; _gv_i_150 = _gv_i_150 + 1) begin : g_execute_out_if
													localparam i = _gv_i_150;
													// Trace: src/VX_pe_switch.sv:41:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[i + _mbase_execute_out_if].valid = pe_req_valid[i];
													// Trace: src/VX_pe_switch.sv:42:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[i + _mbase_execute_out_if].data = pe_req_data[i * 471+:471];
													// Trace: src/VX_pe_switch.sv:43:9
													assign pe_req_ready[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[i + _mbase_execute_out_if].ready;
												end
												// Trace: src/VX_pe_switch.sv:45:5
												wire [1:0] pe_rsp_valid;
												// Trace: src/VX_pe_switch.sv:46:5
												wire [347:0] pe_rsp_data;
												// Trace: src/VX_pe_switch.sv:47:5
												wire [1:0] pe_rsp_ready;
												// Trace: src/VX_pe_switch.sv:48:5
												genvar _gv_i_151;
												for (_gv_i_151 = 0; _gv_i_151 < PE_COUNT; _gv_i_151 = _gv_i_151 + 1) begin : g_result_in_if
													localparam i = _gv_i_151;
													// Trace: src/VX_pe_switch.sv:49:9
													assign pe_rsp_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[i + _mbase_result_in_if].valid;
													// Trace: src/VX_pe_switch.sv:50:9
													assign pe_rsp_data[i * 174+:174] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[i + _mbase_result_in_if].data;
													// Trace: src/VX_pe_switch.sv:51:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[i + _mbase_result_in_if].ready = pe_rsp_ready[i];
												end
												// Trace: src/VX_pe_switch.sv:53:5
												VX_stream_arb #(
													.NUM_INPUTS(PE_COUNT),
													.DATAW(RSP_DATAW),
													.ARBITER(ARBITER),
													.OUT_BUF(RSP_OUT_BUF)
												) rsp_arb(
													.clk(clk),
													.reset(reset),
													.valid_in(pe_rsp_valid),
													.ready_in(pe_rsp_ready),
													.data_in(pe_rsp_data),
													.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_result_if[_mbase_result_out_if].data),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_result_if[_mbase_result_out_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_result_if[_mbase_result_out_if].ready),
													.sel_out()
												);
											end
											assign pe_switch.clk = clk;
											assign pe_switch.reset = reset;
											assign pe_switch.pe_sel = pe_select;
											// Trace: src/VX_alu_unit.sv:61:9
											// expanded module instance: alu_int
											localparam _bbase_EF6D6_execute_if = PE_IDX_INT;
											localparam _bbase_EF6D6_branch_ctl_if = block_idx + _mbase_branch_ctl_if;
											localparam _bbase_EF6D6_result_if = PE_IDX_INT;
											localparam _param_EF6D6_INSTANCE_ID = "";
											localparam _param_EF6D6_BLOCK_IDX = block_idx;
											localparam _param_EF6D6_NUM_LANES = NUM_LANES;
											if (1) begin : alu_int
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_alu_int.sv:2:15
												localparam INSTANCE_ID = _param_EF6D6_INSTANCE_ID;
												// Trace: src/VX_alu_int.sv:3:15
												localparam BLOCK_IDX = _param_EF6D6_BLOCK_IDX;
												// Trace: src/VX_alu_int.sv:4:15
												localparam NUM_LANES = _param_EF6D6_NUM_LANES;
												// Trace: src/VX_alu_int.sv:6:5
												wire clk;
												// Trace: src/VX_alu_int.sv:7:5
												wire reset;
												// Trace: src/VX_alu_int.sv:8:5
												localparam _mbase_execute_if = _bbase_EF6D6_execute_if;
												// Trace: src/VX_alu_int.sv:9:5
												localparam _mbase_result_if = _bbase_EF6D6_result_if;
												// Trace: src/VX_alu_int.sv:10:5
												localparam _mbase_branch_ctl_if = _bbase_EF6D6_branch_ctl_if;
												// Trace: src/VX_alu_int.sv:12:5
												localparam LANE_BITS = 2;
												// Trace: src/VX_alu_int.sv:13:5
												localparam LANE_WIDTH = LANE_BITS;
												// Trace: src/VX_alu_int.sv:14:5
												localparam PID_BITS = 0;
												// Trace: src/VX_alu_int.sv:15:5
												localparam PID_WIDTH = 1;
												// Trace: src/VX_alu_int.sv:16:5
												localparam SHIFT_IMM_BITS = 5;
												// Trace: src/VX_alu_int.sv:17:5
												wire [127:0] add_result;
												// Trace: src/VX_alu_int.sv:18:5
												wire [131:0] sub_result;
												// Trace: src/VX_alu_int.sv:19:5
												reg [127:0] shr_zic_result;
												// Trace: src/VX_alu_int.sv:20:5
												reg [127:0] msc_result;
												// Trace: src/VX_alu_int.sv:21:5
												wire [127:0] add_result_w;
												// Trace: src/VX_alu_int.sv:22:5
												wire [127:0] sub_result_w;
												// Trace: src/VX_alu_int.sv:23:5
												wire [127:0] shr_result_w;
												// Trace: src/VX_alu_int.sv:24:5
												reg [127:0] msc_result_w;
												// Trace: src/VX_alu_int.sv:25:5
												reg [127:0] vote_result;
												// Trace: src/VX_alu_int.sv:26:5
												wire [127:0] shfl_result;
												// Trace: src/VX_alu_int.sv:27:5
												reg [127:0] alu_result;
												// Trace: src/VX_alu_int.sv:28:5
												wire [127:0] alu_result_r;
												// Trace: src/VX_alu_int.sv:29:5
												wire is_alu_w = 0;
												// Trace: src/VX_alu_int.sv:30:5
												localparam VX_gpu_pkg_INST_ALU_BITS = 4;
												wire [3:0] alu_op = sv2v_cast_4(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[433-:4]);
												// Trace: src/VX_alu_int.sv:31:5
												localparam VX_gpu_pkg_INST_BR_BITS = 4;
												wire [3:0] br_op = sv2v_cast_4(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[433-:4]);
												// Trace: src/VX_alu_int.sv:32:5
												localparam VX_gpu_pkg_ALU_TYPE_BRANCH = 1;
												wire is_br_op = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[426-:2] == VX_gpu_pkg_ALU_TYPE_BRANCH;
												// Trace: src/VX_alu_int.sv:33:5
												function automatic VX_gpu_pkg_inst_alu_is_sub;
													// Trace: src/VX_gpu_pkg.sv:120:46
													input reg [3:0] op;
													// Trace: src/VX_gpu_pkg.sv:121:9
													VX_gpu_pkg_inst_alu_is_sub = op[1];
												endfunction
												wire is_sub_op = VX_gpu_pkg_inst_alu_is_sub(alu_op);
												// Trace: src/VX_alu_int.sv:34:5
												function automatic VX_gpu_pkg_inst_alu_signed;
													// Trace: src/VX_gpu_pkg.sv:117:46
													input reg [3:0] op;
													// Trace: src/VX_gpu_pkg.sv:118:9
													VX_gpu_pkg_inst_alu_signed = op[0];
												endfunction
												wire is_signed = VX_gpu_pkg_inst_alu_signed(alu_op);
												// Trace: src/VX_alu_int.sv:35:5
												function automatic [1:0] VX_gpu_pkg_inst_alu_class;
													// Trace: src/VX_gpu_pkg.sv:114:51
													input reg [3:0] op;
													// Trace: src/VX_gpu_pkg.sv:115:9
													VX_gpu_pkg_inst_alu_class = op[3:2];
												endfunction
												function automatic [1:0] VX_gpu_pkg_inst_br_class;
													// Trace: src/VX_gpu_pkg.sv:141:50
													input reg [3:0] op;
													// Trace: src/VX_gpu_pkg.sv:142:9
													VX_gpu_pkg_inst_br_class = {1'b0, ~op[3]};
												endfunction
												wire [1:0] op_class = (is_br_op ? VX_gpu_pkg_inst_br_class(alu_op) : VX_gpu_pkg_inst_alu_class(alu_op));
												// Trace: src/VX_alu_int.sv:36:5
												wire [127:0] alu_in1 = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[386-:128];
												// Trace: src/VX_alu_int.sv:37:5
												wire [127:0] alu_in2 = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[258-:128];
												// Trace: src/VX_alu_int.sv:38:5
												localparam VX_gpu_pkg_PC_BITS = 30;
												function automatic [31:0] VX_gpu_pkg_to_fullPC;
													// Trace: src/VX_gpu_pkg.sv:27:49
													input reg [29:0] pc;
													// Trace: src/VX_gpu_pkg.sv:28:9
													VX_gpu_pkg_to_fullPC = {pc, 2'b00};
												endfunction
												wire [127:0] alu_in1_PC = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[429] ? {NUM_LANES {VX_gpu_pkg_to_fullPC(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[463-:30])}} : alu_in1);
												// Trace: src/VX_alu_int.sv:39:5
												wire [127:0] alu_in2_imm = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[428] ? {NUM_LANES {{Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[424], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[423:393]}}} : alu_in2);
												// Trace: src/VX_alu_int.sv:40:5
												wire [127:0] alu_in2_br = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[428] && ~is_br_op ? {NUM_LANES {{Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[424], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[423:393]}}} : alu_in2);
												// Trace: src/VX_alu_int.sv:41:5
												genvar _gv_i_141;
												for (_gv_i_141 = 0; _gv_i_141 < NUM_LANES; _gv_i_141 = _gv_i_141 + 1) begin : g_add_result
													localparam i = _gv_i_141;
													// Trace: src/VX_alu_int.sv:42:9
													assign add_result[i * 32+:32] = alu_in1_PC[i * 32+:32] + alu_in2_imm[i * 32+:32];
													// Trace: src/VX_alu_int.sv:43:9
													assign add_result_w[i * 32+:32] = sv2v_cast_32_signed($signed(alu_in1[(i * 32) + 31-:32] + alu_in2_imm[(i * 32) + 31-:32]));
												end
												// Trace: src/VX_alu_int.sv:45:5
												genvar _gv_i_142;
												for (_gv_i_142 = 0; _gv_i_142 < NUM_LANES; _gv_i_142 = _gv_i_142 + 1) begin : g_sub_result
													localparam i = _gv_i_142;
													// Trace: src/VX_alu_int.sv:46:9
													wire [32:0] sub_in1 = {is_signed & alu_in1[(i * 32) + 31], alu_in1[i * 32+:32]};
													// Trace: src/VX_alu_int.sv:47:9
													wire [32:0] sub_in2 = {is_signed & alu_in2_br[(i * 32) + 31], alu_in2_br[i * 32+:32]};
													// Trace: src/VX_alu_int.sv:48:9
													assign sub_result[i * 33+:33] = sub_in1 - sub_in2;
													// Trace: src/VX_alu_int.sv:49:9
													assign sub_result_w[i * 32+:32] = sv2v_cast_32_signed($signed(alu_in1[(i * 32) + 31-:32] - alu_in2_imm[(i * 32) + 31-:32]));
												end
												// Trace: src/VX_alu_int.sv:51:5
												genvar _gv_i_143;
												for (_gv_i_143 = 0; _gv_i_143 < NUM_LANES; _gv_i_143 = _gv_i_143 + 1) begin : g_shr_result
													localparam i = _gv_i_143;
													// Trace: src/VX_alu_int.sv:52:9
													wire [32:0] shr_in1 = {is_signed && alu_in1[(i * 32) + 31], alu_in1[i * 32+:32]};
													// Trace: src/VX_alu_int.sv:53:9
													always @(*)
														// Trace: src/VX_alu_int.sv:54:13
														case (alu_op[1:0])
															2'b10, 2'b11:
																// Trace: src/VX_alu_int.sv:56:21
																shr_zic_result[i * 32+:32] = alu_in1[i * 32+:32] & {32 {alu_op[0] ^ |alu_in2[i * 32+:32]}};
															default:
																// Trace: src/VX_alu_int.sv:59:21
																shr_zic_result[i * 32+:32] = sv2v_cast_32_signed($signed(shr_in1) >>> alu_in2_imm[(i * 32) + 4-:5]);
														endcase
													// Trace: src/VX_alu_int.sv:63:9
													wire [32:0] shr_in1_w = {is_signed && alu_in1[(i * 32) + 31], alu_in1[(i * 32) + 31-:32]};
													// Trace: src/VX_alu_int.sv:64:9
													wire [31:0] shr_res_w = sv2v_cast_32_signed($signed(shr_in1_w) >>> alu_in2_imm[(i * 32) + 4-:5]);
													// Trace: src/VX_alu_int.sv:65:9
													assign shr_result_w[i * 32+:32] = sv2v_cast_32_signed($signed(shr_res_w));
												end
												// Trace: src/VX_alu_int.sv:67:5
												genvar _gv_i_144;
												for (_gv_i_144 = 0; _gv_i_144 < NUM_LANES; _gv_i_144 = _gv_i_144 + 1) begin : g_msc_result
													localparam i = _gv_i_144;
													// Trace: src/VX_alu_int.sv:68:9
													always @(*)
														// Trace: src/VX_alu_int.sv:69:13
														case (alu_op[1:0])
															2'b00:
																// Trace: src/VX_alu_int.sv:70:24
																msc_result[i * 32+:32] = alu_in1[i * 32+:32] & alu_in2_imm[i * 32+:32];
															2'b01:
																// Trace: src/VX_alu_int.sv:71:24
																msc_result[i * 32+:32] = alu_in1[i * 32+:32] | alu_in2_imm[i * 32+:32];
															2'b10:
																// Trace: src/VX_alu_int.sv:72:24
																msc_result[i * 32+:32] = alu_in1[i * 32+:32] ^ alu_in2_imm[i * 32+:32];
															2'b11:
																// Trace: src/VX_alu_int.sv:73:24
																msc_result[i * 32+:32] = alu_in1[i * 32+:32] << alu_in2_imm[(i * 32) + 4-:5];
														endcase
													// Trace: src/VX_alu_int.sv:76:9
													wire [32:1] sv2v_tmp_4E506;
													assign sv2v_tmp_4E506 = sv2v_cast_32_signed($signed(alu_in1[(i * 32) + 31-:32] << alu_in2_imm[(i * 32) + 4-:5]));
													always @(*) msc_result_w[i * 32+:32] = sv2v_tmp_4E506;
												end
												// Trace: src/VX_alu_int.sv:78:5
												wire [3:0] vote_true;
												wire [3:0] vote_false;
												// Trace: src/VX_alu_int.sv:79:5
												genvar _gv_i_145;
												for (_gv_i_145 = 0; _gv_i_145 < NUM_LANES; _gv_i_145 = _gv_i_145 + 1) begin : g_vote_calc
													localparam i = _gv_i_145;
													// Trace: src/VX_alu_int.sv:80:9
													wire pred = alu_in1[i * 32];
													// Trace: src/VX_alu_int.sv:81:9
													assign vote_true[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[464 + i] && pred;
													// Trace: src/VX_alu_int.sv:82:9
													assign vote_false[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[464 + i] && ~pred;
												end
												// Trace: src/VX_alu_int.sv:84:5
												wire has_vote_true = |vote_true;
												// Trace: src/VX_alu_int.sv:85:5
												wire has_vote_false = |vote_false;
												// Trace: src/VX_alu_int.sv:86:5
												wire vote_all = ~has_vote_false;
												// Trace: src/VX_alu_int.sv:87:5
												wire vote_any = has_vote_true;
												// Trace: src/VX_alu_int.sv:88:5
												wire vote_none = ~has_vote_true;
												// Trace: src/VX_alu_int.sv:89:5
												wire vote_uni = vote_all || vote_none;
												// Trace: src/VX_alu_int.sv:90:5
												genvar _gv_i_146;
												localparam VX_gpu_pkg_INST_VOTE_ALL = 2'b00;
												localparam VX_gpu_pkg_INST_VOTE_ANY = 2'b01;
												localparam VX_gpu_pkg_INST_VOTE_BAL = 2'b11;
												localparam VX_gpu_pkg_INST_VOTE_UNI = 2'b10;
												for (_gv_i_146 = 0; _gv_i_146 < NUM_LANES; _gv_i_146 = _gv_i_146 + 1) begin : g_vote_result
													localparam i = _gv_i_146;
													// Trace: src/VX_alu_int.sv:91:9
													always @(*)
														// Trace: src/VX_alu_int.sv:92:13
														case (alu_op[1:0])
															VX_gpu_pkg_INST_VOTE_ALL:
																// Trace: src/VX_alu_int.sv:93:32
																vote_result[i * 32+:32] = sv2v_cast_32(vote_all);
															VX_gpu_pkg_INST_VOTE_ANY:
																// Trace: src/VX_alu_int.sv:94:32
																vote_result[i * 32+:32] = sv2v_cast_32(vote_any);
															VX_gpu_pkg_INST_VOTE_UNI:
																// Trace: src/VX_alu_int.sv:95:32
																vote_result[i * 32+:32] = sv2v_cast_32(vote_uni);
															VX_gpu_pkg_INST_VOTE_BAL:
																// Trace: src/VX_alu_int.sv:96:32
																vote_result[i * 32+:32] = sv2v_cast_32(vote_true);
														endcase
												end
												// Trace: src/VX_alu_int.sv:100:5
												localparam VX_gpu_pkg_INST_SHFL_BFLY = 2'b10;
												localparam VX_gpu_pkg_INST_SHFL_DOWN = 2'b01;
												localparam VX_gpu_pkg_INST_SHFL_IDX = 2'b11;
												localparam VX_gpu_pkg_INST_SHFL_UP = 2'b00;
												if (1) begin : g_shfl
													genvar _gv_i_147;
													for (_gv_i_147 = 0; _gv_i_147 < NUM_LANES; _gv_i_147 = _gv_i_147 + 1) begin : g_i
														localparam i = _gv_i_147;
														// Trace: src/VX_alu_int.sv:102:13
														wire [1:0] bval = alu_in2[i * 32+:LANE_BITS];
														// Trace: src/VX_alu_int.sv:103:13
														wire [1:0] cval = alu_in2[(i * 32) + 6+:LANE_BITS];
														// Trace: src/VX_alu_int.sv:104:13
														wire [1:0] mask = alu_in2[(i * 32) + 12+:LANE_BITS];
														// Trace: src/VX_alu_int.sv:105:13
														wire [1:0] minLane = sv2v_cast_2_signed(i) & mask;
														// Trace: src/VX_alu_int.sv:106:13
														wire [1:0] maxLane = minLane | (cval & ~mask);
														// Trace: src/VX_alu_int.sv:107:13
														wire [LANE_BITS:0] lane_up = sv2v_cast_2_signed(i) - bval;
														// Trace: src/VX_alu_int.sv:108:13
														wire [LANE_BITS:0] lane_down = sv2v_cast_2_signed(i) + bval;
														// Trace: src/VX_alu_int.sv:109:13
														wire [1:0] lane_bfly = sv2v_cast_2_signed(i) ^ bval;
														// Trace: src/VX_alu_int.sv:110:13
														wire [1:0] lane_idx = minLane | (bval & ~mask);
														// Trace: src/VX_alu_int.sv:111:13
														reg [1:0] lane;
														// Trace: src/VX_alu_int.sv:112:13
														always @(*) begin
															// Trace: src/VX_alu_int.sv:113:17
															lane = sv2v_cast_2_signed(i);
															// Trace: src/VX_alu_int.sv:114:17
															case (alu_op[1:0])
																VX_gpu_pkg_INST_SHFL_UP:
																	// Trace: src/VX_alu_int.sv:116:25
																	if ($signed(lane_up) >= $signed({1'b0, minLane}))
																		// Trace: src/VX_alu_int.sv:117:29
																		lane = lane_up[1:0];
																VX_gpu_pkg_INST_SHFL_DOWN:
																	// Trace: src/VX_alu_int.sv:121:25
																	if (lane_down <= {1'b0, maxLane})
																		// Trace: src/VX_alu_int.sv:122:29
																		lane = lane_down[1:0];
																VX_gpu_pkg_INST_SHFL_BFLY:
																	// Trace: src/VX_alu_int.sv:126:25
																	if (lane_bfly <= maxLane)
																		// Trace: src/VX_alu_int.sv:127:29
																		lane = lane_bfly;
																VX_gpu_pkg_INST_SHFL_IDX:
																	// Trace: src/VX_alu_int.sv:131:25
																	if (lane_idx <= maxLane)
																		// Trace: src/VX_alu_int.sv:132:29
																		lane = lane_idx;
															endcase
														end
														// Trace: src/VX_alu_int.sv:137:13
														assign shfl_result[i * 32+:32] = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[0].data[464 + lane] ? alu_in1[lane * 32+:32] : alu_in1[i * 32+:32]);
													end
												end
												// Trace: src/VX_alu_int.sv:142:5
												genvar _gv_i_148;
												localparam VX_gpu_pkg_ALU_TYPE_OTHER = 3;
												for (_gv_i_148 = 0; _gv_i_148 < NUM_LANES; _gv_i_148 = _gv_i_148 + 1) begin : g_alu_result
													localparam i = _gv_i_148;
													// Trace: src/VX_alu_int.sv:143:9
													wire [31:0] slt_br_result = sv2v_cast_32({is_br_op && ~(|sub_result[(i * 33) + 31-:32]), sub_result[(i * 33) + 32]});
													// Trace: src/VX_alu_int.sv:144:9
													wire [31:0] sub_slt_br_result = (is_sub_op && ~is_br_op ? sub_result[(i * 33) + 31-:32] : slt_br_result);
													// Trace: src/VX_alu_int.sv:145:9
													always @(*)
														// Trace: src/VX_alu_int.sv:146:13
														if (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[426-:2] == VX_gpu_pkg_ALU_TYPE_OTHER)
															// Trace: src/VX_alu_int.sv:147:17
															case (alu_op[2])
																1'b0:
																	// Trace: src/VX_alu_int.sv:148:27
																	alu_result[i * 32+:32] = vote_result[i * 32+:32];
																1'b1:
																	// Trace: src/VX_alu_int.sv:149:27
																	alu_result[i * 32+:32] = shfl_result[i * 32+:32];
																default:
																	;
															endcase
														else
															// Trace: src/VX_alu_int.sv:153:17
															case ({is_alu_w, op_class})
																3'b000:
																	// Trace: src/VX_alu_int.sv:154:29
																	alu_result[i * 32+:32] = add_result[i * 32+:32];
																3'b001:
																	// Trace: src/VX_alu_int.sv:155:29
																	alu_result[i * 32+:32] = sub_slt_br_result;
																3'b010:
																	// Trace: src/VX_alu_int.sv:156:29
																	alu_result[i * 32+:32] = shr_zic_result[i * 32+:32];
																3'b011:
																	// Trace: src/VX_alu_int.sv:157:29
																	alu_result[i * 32+:32] = msc_result[i * 32+:32];
																3'b100:
																	// Trace: src/VX_alu_int.sv:158:29
																	alu_result[i * 32+:32] = add_result_w[i * 32+:32];
																3'b101:
																	// Trace: src/VX_alu_int.sv:159:29
																	alu_result[i * 32+:32] = sub_result_w[i * 32+:32];
																3'b110:
																	// Trace: src/VX_alu_int.sv:160:29
																	alu_result[i * 32+:32] = shr_result_w[i * 32+:32];
																3'b111:
																	// Trace: src/VX_alu_int.sv:161:29
																	alu_result[i * 32+:32] = msc_result_w[i * 32+:32];
															endcase
												end
												// Trace: src/VX_alu_int.sv:166:5
												wire [29:0] PC_r;
												// Trace: src/VX_alu_int.sv:167:5
												wire [3:0] br_op_r;
												// Trace: src/VX_alu_int.sv:168:5
												wire [29:0] cbr_dest;
												wire [29:0] cbr_dest_r;
												// Trace: src/VX_alu_int.sv:169:5
												wire [1:0] last_tid;
												wire [1:0] last_tid_r;
												// Trace: src/VX_alu_int.sv:170:5
												wire is_br_op_r;
												// Trace: src/VX_alu_int.sv:171:5
												function automatic [29:0] VX_gpu_pkg_from_fullPC;
													// Trace: src/VX_gpu_pkg.sv:30:56
													input reg [31:0] pc;
													// Trace: src/VX_gpu_pkg.sv:31:9
													VX_gpu_pkg_from_fullPC = sv2v_cast_30(pc >> 2);
												endfunction
												assign cbr_dest = VX_gpu_pkg_from_fullPC(add_result[0+:32]);
												// Trace: src/VX_alu_int.sv:172:5
												if (1) begin : g_last_tid
													// Trace: src/VX_alu_int.sv:173:9
													VX_priority_encoder #(
														.N(NUM_LANES),
														.REVERSE(1)
													) last_tid_sel(
														.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[467-:4]),
														.index_out(last_tid),
														.onehot_out(),
														.valid_out()
													);
												end
												// Trace: src/VX_alu_int.sv:185:5
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_RV_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
												localparam VX_gpu_pkg_NW_BITS = 2;
												localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												VX_elastic_buffer #(.DATAW(211)) rsp_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].valid),
													.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].ready),
													.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[470], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[469-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[467-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[391-:5], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[392], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[0], alu_result, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[463-:30], cbr_dest, is_br_op, br_op, last_tid}),
													.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[173], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[172-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[170-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[135-:5], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[136], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[0], alu_result_r, PC_r, cbr_dest_r, is_br_op_r, br_op_r, last_tid_r}),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].ready)
												);
												// Trace: src/VX_alu_int.sv:197:5
												function automatic VX_gpu_pkg_inst_br_is_neg;
													// Trace: src/VX_gpu_pkg.sv:144:45
													input reg [3:0] op;
													// Trace: src/VX_gpu_pkg.sv:145:9
													VX_gpu_pkg_inst_br_is_neg = op[1];
												endfunction
												wire is_br_neg = VX_gpu_pkg_inst_br_is_neg(br_op_r);
												// Trace: src/VX_alu_int.sv:198:5
												function automatic VX_gpu_pkg_inst_br_is_less;
													// Trace: src/VX_gpu_pkg.sv:147:46
													input reg [3:0] op;
													// Trace: src/VX_gpu_pkg.sv:148:9
													VX_gpu_pkg_inst_br_is_less = op[2];
												endfunction
												wire is_br_less = VX_gpu_pkg_inst_br_is_less(br_op_r);
												// Trace: src/VX_alu_int.sv:199:5
												function automatic VX_gpu_pkg_inst_br_is_static;
													// Trace: src/VX_gpu_pkg.sv:150:48
													input reg [3:0] op;
													// Trace: src/VX_gpu_pkg.sv:151:9
													VX_gpu_pkg_inst_br_is_static = op[3];
												endfunction
												wire is_br_static = VX_gpu_pkg_inst_br_is_static(br_op_r);
												// Trace: src/VX_alu_int.sv:200:5
												wire [31:0] br_result = alu_result_r[last_tid_r * 32+:32];
												// Trace: src/VX_alu_int.sv:201:5
												wire is_less = br_result[0];
												// Trace: src/VX_alu_int.sv:202:5
												wire is_equal = br_result[1];
												// Trace: src/VX_alu_int.sv:203:5
												wire result_fire = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].ready;
												// Trace: src/VX_alu_int.sv:204:5
												wire br_enable = (result_fire && is_br_op_r) && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[0];
												// Trace: src/VX_alu_int.sv:205:5
												wire br_taken = ((is_br_less ? is_less : is_equal) ^ is_br_neg) | is_br_static;
												// Trace: src/VX_alu_int.sv:206:5
												wire [29:0] br_dest = (is_br_static ? VX_gpu_pkg_from_fullPC(br_result) : cbr_dest_r);
												// Trace: src/VX_alu_int.sv:207:5
												wire [1:0] br_wid;
												// Trace: src/VX_alu_int.sv:209:5
												if (1) begin : genblk10
													// Trace: src/VX_alu_int.sv:216:9
													assign br_wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[172-:2];
												end
												// Trace: src/VX_alu_int.sv:219:5
												VX_pipe_register #(
													.DATAW(34),
													.RESETW(1)
												) branch_reg(
													.clk(clk),
													.reset(reset),
													.enable(1'b1),
													.data_in({br_enable, br_wid, br_taken, br_dest}),
													.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[_mbase_branch_ctl_if].valid, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[_mbase_branch_ctl_if].wid, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[_mbase_branch_ctl_if].taken, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.branch_ctl_if[_mbase_branch_ctl_if].dest})
												);
												// Trace: src/VX_alu_int.sv:229:5
												genvar _gv_i_149;
												for (_gv_i_149 = 0; _gv_i_149 < NUM_LANES; _gv_i_149 = _gv_i_149 + 1) begin : g_result
													localparam i = _gv_i_149;
													// Trace: src/VX_alu_int.sv:230:9
													wire [31:0] PC_next = VX_gpu_pkg_to_fullPC(PC_r) + 32'sd4;
													// Trace: src/VX_alu_int.sv:231:9
													assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[3 + (i * 32)+:32] = (is_br_op_r && is_br_static ? PC_next : alu_result_r[i * 32+:32]);
												end
												// Trace: src/VX_alu_int.sv:233:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[166-:30] = PC_r;
											end
											assign alu_int.clk = clk;
											assign alu_int.reset = reset;
											// Trace: src/VX_alu_unit.sv:72:9
											// expanded module instance: muldiv_unit
											localparam _bbase_50917_execute_if = PE_IDX_MDV;
											localparam _bbase_50917_result_if = PE_IDX_MDV;
											localparam _param_50917_INSTANCE_ID = "";
											localparam _param_50917_NUM_LANES = NUM_LANES;
											if (1) begin : muldiv_unit
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_alu_muldiv.sv:2:15
												localparam INSTANCE_ID = _param_50917_INSTANCE_ID;
												// Trace: src/VX_alu_muldiv.sv:3:15
												localparam NUM_LANES = _param_50917_NUM_LANES;
												// Trace: src/VX_alu_muldiv.sv:5:5
												wire clk;
												// Trace: src/VX_alu_muldiv.sv:6:5
												wire reset;
												// Trace: src/VX_alu_muldiv.sv:7:5
												localparam _mbase_execute_if = _bbase_50917_execute_if;
												// Trace: src/VX_alu_muldiv.sv:8:5
												localparam _mbase_result_if = _bbase_50917_result_if;
												// Trace: src/VX_alu_muldiv.sv:10:5
												localparam PID_BITS = 0;
												// Trace: src/VX_alu_muldiv.sv:11:5
												localparam PID_WIDTH = 1;
												// Trace: src/VX_alu_muldiv.sv:12:5
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_RV_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
												localparam VX_gpu_pkg_NW_BITS = 2;
												localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
												localparam VX_gpu_pkg_PC_BITS = 30;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam TAG_WIDTH = 46;
												// Trace: src/VX_alu_muldiv.sv:13:5
												localparam VX_gpu_pkg_INST_M_BITS = 3;
												wire [2:0] muldiv_op = sv2v_cast_3(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[433-:4]);
												// Trace: src/VX_alu_muldiv.sv:14:5
												function automatic VX_gpu_pkg_inst_m_is_mulx;
													// Trace: src/VX_gpu_pkg.sv:175:45
													input reg [2:0] op;
													// Trace: src/VX_gpu_pkg.sv:176:9
													VX_gpu_pkg_inst_m_is_mulx = ~op[2];
												endfunction
												wire is_mulx_op = VX_gpu_pkg_inst_m_is_mulx(muldiv_op);
												// Trace: src/VX_alu_muldiv.sv:15:5
												function automatic VX_gpu_pkg_inst_m_signed;
													// Trace: src/VX_gpu_pkg.sv:172:44
													input reg [2:0] op;
													// Trace: src/VX_gpu_pkg.sv:173:9
													VX_gpu_pkg_inst_m_signed = ~op[0];
												endfunction
												wire is_signed_op = VX_gpu_pkg_inst_m_signed(muldiv_op);
												// Trace: src/VX_alu_muldiv.sv:16:5
												wire is_alu_w = 0;
												// Trace: src/VX_alu_muldiv.sv:17:5
												wire [127:0] mul_result_out;
												// Trace: src/VX_alu_muldiv.sv:18:5
												wire [0:0] mul_uuid_out;
												// Trace: src/VX_alu_muldiv.sv:19:5
												wire [1:0] mul_wid_out;
												// Trace: src/VX_alu_muldiv.sv:20:5
												wire [3:0] mul_tmask_out;
												// Trace: src/VX_alu_muldiv.sv:21:5
												wire [29:0] mul_PC_out;
												// Trace: src/VX_alu_muldiv.sv:22:5
												wire [4:0] mul_rd_out;
												// Trace: src/VX_alu_muldiv.sv:23:5
												wire mul_wb_out;
												// Trace: src/VX_alu_muldiv.sv:24:5
												wire [0:0] mul_pid_out;
												// Trace: src/VX_alu_muldiv.sv:25:5
												wire mul_sop_out;
												wire mul_eop_out;
												// Trace: src/VX_alu_muldiv.sv:26:5
												wire mul_valid_in = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].valid && is_mulx_op;
												// Trace: src/VX_alu_muldiv.sv:27:5
												wire mul_ready_in;
												// Trace: src/VX_alu_muldiv.sv:28:5
												wire mul_valid_out;
												// Trace: src/VX_alu_muldiv.sv:29:5
												wire mul_ready_out;
												// Trace: src/VX_alu_muldiv.sv:30:5
												function automatic VX_gpu_pkg_inst_m_is_mulh;
													// Trace: src/VX_gpu_pkg.sv:178:45
													input reg [2:0] op;
													// Trace: src/VX_gpu_pkg.sv:179:9
													VX_gpu_pkg_inst_m_is_mulh = op[1:0] != 0;
												endfunction
												wire is_mulh_in = VX_gpu_pkg_inst_m_is_mulh(muldiv_op);
												// Trace: src/VX_alu_muldiv.sv:31:5
												function automatic VX_gpu_pkg_inst_m_signed_a;
													// Trace: src/VX_gpu_pkg.sv:181:46
													input reg [2:0] op;
													// Trace: src/VX_gpu_pkg.sv:182:9
													VX_gpu_pkg_inst_m_signed_a = op[1:0] != 1;
												endfunction
												wire is_signed_mul_a = VX_gpu_pkg_inst_m_signed_a(muldiv_op);
												// Trace: src/VX_alu_muldiv.sv:32:5
												wire is_signed_mul_b = is_signed_op;
												// Trace: src/VX_alu_muldiv.sv:33:5
												wire [263:0] mul_result_tmp;
												// Trace: src/VX_alu_muldiv.sv:34:5
												wire is_mulh_out;
												// Trace: src/VX_alu_muldiv.sv:35:5
												wire is_mul_w_out;
												// Trace: src/VX_alu_muldiv.sv:36:5
												genvar _gv_i_76;
												for (_gv_i_76 = 0; _gv_i_76 < NUM_LANES; _gv_i_76 = _gv_i_76 + 1) begin : g_multiplier
													localparam i = _gv_i_76;
													// Trace: src/VX_alu_muldiv.sv:37:9
													wire [32:0] mul_in1 = {is_signed_mul_a && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[259 + ((i * 32) + 31)], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[259 + (i * 32)+:32]};
													// Trace: src/VX_alu_muldiv.sv:38:9
													wire [32:0] mul_in2 = {is_signed_mul_b && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[131 + ((i * 32) + 31)], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[131 + (i * 32)+:32]};
													// Trace: src/VX_alu_muldiv.sv:39:9
													VX_multiplier #(
														.A_WIDTH(33),
														.B_WIDTH(33),
														.R_WIDTH(66),
														.SIGNED(1),
														.LATENCY(3)
													) multiplier(
														.clk(clk),
														.enable(mul_ready_in),
														.dataa(mul_in1),
														.datab(mul_in2),
														.result(mul_result_tmp[i * 66+:66])
													);
												end
												// Trace: src/VX_alu_muldiv.sv:53:5
												VX_shift_register #(
													.DATAW(49),
													.DEPTH(3),
													.RESETW(1)
												) mul_shift_reg(
													.clk(clk),
													.reset(reset),
													.enable(mul_ready_in),
													.data_in({mul_valid_in, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[470], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[469-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[467-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[463-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[391-:5], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[392], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[0], is_mulh_in, is_alu_w}),
													.data_out({mul_valid_out, mul_uuid_out, mul_wid_out, mul_tmask_out, mul_PC_out, mul_rd_out, mul_wb_out, mul_pid_out, mul_sop_out, mul_eop_out, is_mulh_out, is_mul_w_out})
												);
												// Trace: src/VX_alu_muldiv.sv:64:5
												assign mul_ready_in = mul_ready_out || ~mul_valid_out;
												// Trace: src/VX_alu_muldiv.sv:65:5
												genvar _gv_i_77;
												for (_gv_i_77 = 0; _gv_i_77 < NUM_LANES; _gv_i_77 = _gv_i_77 + 1) begin : g_mul_result_out
													localparam i = _gv_i_77;
													// Trace: src/VX_alu_muldiv.sv:66:9
													assign mul_result_out[i * 32+:32] = (is_mulh_out ? mul_result_tmp[(i * 66) + 63-:32] : mul_result_tmp[(i * 66) + 31-:32]);
												end
												// Trace: src/VX_alu_muldiv.sv:68:5
												wire [127:0] div_result_out;
												// Trace: src/VX_alu_muldiv.sv:69:5
												wire [0:0] div_uuid_out;
												// Trace: src/VX_alu_muldiv.sv:70:5
												wire [1:0] div_wid_out;
												// Trace: src/VX_alu_muldiv.sv:71:5
												wire [3:0] div_tmask_out;
												// Trace: src/VX_alu_muldiv.sv:72:5
												wire [29:0] div_PC_out;
												// Trace: src/VX_alu_muldiv.sv:73:5
												wire [4:0] div_rd_out;
												// Trace: src/VX_alu_muldiv.sv:74:5
												wire div_wb_out;
												// Trace: src/VX_alu_muldiv.sv:75:5
												wire [0:0] div_pid_out;
												// Trace: src/VX_alu_muldiv.sv:76:5
												wire div_sop_out;
												wire div_eop_out;
												// Trace: src/VX_alu_muldiv.sv:77:5
												function automatic VX_gpu_pkg_inst_m_is_rem;
													// Trace: src/VX_gpu_pkg.sv:184:44
													input reg [2:0] op;
													// Trace: src/VX_gpu_pkg.sv:185:9
													VX_gpu_pkg_inst_m_is_rem = op[1];
												endfunction
												wire is_rem_op = VX_gpu_pkg_inst_m_is_rem(muldiv_op);
												// Trace: src/VX_alu_muldiv.sv:78:5
												wire div_valid_in = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].valid && ~is_mulx_op;
												// Trace: src/VX_alu_muldiv.sv:79:5
												wire div_ready_in;
												// Trace: src/VX_alu_muldiv.sv:80:5
												wire div_valid_out;
												// Trace: src/VX_alu_muldiv.sv:81:5
												wire div_ready_out;
												// Trace: src/VX_alu_muldiv.sv:82:5
												wire [127:0] div_in1;
												// Trace: src/VX_alu_muldiv.sv:83:5
												wire [127:0] div_in2;
												// Trace: src/VX_alu_muldiv.sv:84:5
												genvar _gv_i_78;
												for (_gv_i_78 = 0; _gv_i_78 < NUM_LANES; _gv_i_78 = _gv_i_78 + 1) begin : g_div_in
													localparam i = _gv_i_78;
													// Trace: src/VX_alu_muldiv.sv:85:9
													assign div_in1[i * 32+:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[259 + (i * 32)+:32];
													// Trace: src/VX_alu_muldiv.sv:86:9
													assign div_in2[i * 32+:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[131 + (i * 32)+:32];
												end
												// Trace: src/VX_alu_muldiv.sv:88:5
												wire [127:0] div_quotient;
												wire [127:0] div_remainder;
												// Trace: src/VX_alu_muldiv.sv:89:5
												wire is_rem_op_out;
												// Trace: src/VX_alu_muldiv.sv:90:5
												wire is_div_w_out;
												// Trace: src/VX_alu_muldiv.sv:91:5
												wire div_strode;
												// Trace: src/VX_alu_muldiv.sv:92:5
												wire div_busy;
												// Trace: src/VX_alu_muldiv.sv:93:5
												VX_elastic_adapter div_elastic_adapter(
													.clk(clk),
													.reset(reset),
													.valid_in(div_valid_in),
													.ready_in(div_ready_in),
													.valid_out(div_valid_out),
													.ready_out(div_ready_out),
													.strobe(div_strode),
													.busy(div_busy)
												);
												// Trace: src/VX_alu_muldiv.sv:103:5
												VX_serial_div #(
													.WIDTHN(32),
													.WIDTHD(32),
													.WIDTHQ(32),
													.WIDTHR(32),
													.LANES(NUM_LANES)
												) serial_div(
													.clk(clk),
													.reset(reset),
													.strobe(div_strode),
													.busy(div_busy),
													.is_signed(is_signed_op),
													.numer(div_in1),
													.denom(div_in2),
													.quotient(div_quotient),
													.remainder(div_remainder)
												);
												// Trace: src/VX_alu_muldiv.sv:120:5
												reg [47:0] div_tag_r;
												// Trace: src/VX_alu_muldiv.sv:121:5
												always @(posedge clk)
													// Trace: src/VX_alu_muldiv.sv:122:9
													if (div_valid_in && div_ready_in)
														// Trace: src/VX_alu_muldiv.sv:123:13
														div_tag_r <= {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[470], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[469-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[467-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[463-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[391-:5], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[392], is_rem_op, is_alu_w, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].data[0]};
												// Trace: src/VX_alu_muldiv.sv:126:5
												assign {div_uuid_out, div_wid_out, div_tmask_out, div_PC_out, div_rd_out, div_wb_out, is_rem_op_out, is_div_w_out, div_pid_out, div_sop_out, div_eop_out} = div_tag_r;
												// Trace: src/VX_alu_muldiv.sv:127:5
												genvar _gv_i_79;
												for (_gv_i_79 = 0; _gv_i_79 < NUM_LANES; _gv_i_79 = _gv_i_79 + 1) begin : g_div_result_out
													localparam i = _gv_i_79;
													// Trace: src/VX_alu_muldiv.sv:128:9
													assign div_result_out[i * 32+:32] = (is_rem_op_out ? div_remainder[i * 32+:32] : div_quotient[i * 32+:32]);
												end
												// Trace: src/VX_alu_muldiv.sv:130:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_execute_if[_mbase_execute_if].ready = (is_mulx_op ? mul_ready_in : div_ready_in);
												// Trace: src/VX_alu_muldiv.sv:131:5
												VX_stream_arb #(
													.NUM_INPUTS(2),
													.DATAW(174),
													.ARBITER("P"),
													.OUT_BUF(2)
												) rsp_buf(
													.clk(clk),
													.reset(reset),
													.valid_in({div_valid_out, mul_valid_out}),
													.ready_in({div_ready_out, mul_ready_out}),
													.data_in({div_uuid_out, div_wid_out, div_tmask_out, div_PC_out, div_rd_out, div_wb_out, div_pid_out, div_sop_out, div_eop_out, div_result_out, mul_uuid_out, mul_wid_out, mul_tmask_out, mul_PC_out, mul_rd_out, mul_wb_out, mul_pid_out, mul_sop_out, mul_eop_out, mul_result_out}),
													.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[173], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[172-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[170-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[166-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[135-:5], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[136], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[0], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].data[130-:128]}),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.g_blocks[_gv_block_idx_1].pe_result_if[_mbase_result_if].ready),
													.sel_out()
												);
											end
											assign muldiv_unit.clk = clk;
											assign muldiv_unit.reset = reset;
										end
										// Trace: src/VX_alu_unit.sv:82:5
										// expanded module instance: gather_unit
										localparam _bbase_8E516_result_if = 0;
										localparam _bbase_8E516_commit_if = 0;
										localparam _param_8E516_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_8E516_NUM_LANES = NUM_LANES;
										localparam _param_8E516_OUT_BUF = (PARTIAL_BW ? 3 : 0);
										if (1) begin : gather_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_gather_unit.sv:2:15
											localparam BLOCK_SIZE = _param_8E516_BLOCK_SIZE;
											// Trace: src/VX_gather_unit.sv:3:15
											localparam NUM_LANES = _param_8E516_NUM_LANES;
											// Trace: src/VX_gather_unit.sv:4:15
											localparam OUT_BUF = _param_8E516_OUT_BUF;
											// Trace: src/VX_gather_unit.sv:6:5
											wire clk;
											// Trace: src/VX_gather_unit.sv:7:5
											wire reset;
											// Trace: src/VX_gather_unit.sv:8:5
											localparam _mbase_result_if = 0;
											// Trace: src/VX_gather_unit.sv:9:5
											localparam _mbase_commit_if = 0;
											// Trace: src/VX_gather_unit.sv:11:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_gather_unit.sv:12:5
											localparam NUM_PACKETS = 1;
											// Trace: src/VX_gather_unit.sv:13:5
											localparam LPID_BITS = 0;
											// Trace: src/VX_gather_unit.sv:14:5
											localparam LPID_WIDTH = 1;
											// Trace: src/VX_gather_unit.sv:15:5
											localparam GPID_BITS = 0;
											// Trace: src/VX_gather_unit.sv:16:5
											localparam GPID_WIDTH = 1;
											// Trace: src/VX_gather_unit.sv:17:5
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam DATAW = 174;
											// Trace: src/VX_gather_unit.sv:18:5
											localparam DATA_WIS_OFF = 171;
											// Trace: src/VX_gather_unit.sv:19:5
											wire [0:0] result_in_valid;
											// Trace: src/VX_gather_unit.sv:20:5
											wire [173:0] result_in_data;
											// Trace: src/VX_gather_unit.sv:21:5
											wire [0:0] result_in_ready;
											// Trace: src/VX_gather_unit.sv:22:5
											localparam VX_gpu_pkg_ISSUE_ISW_BITS = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											wire [0:0] result_in_isw;
											// Trace: src/VX_gather_unit.sv:23:5
											genvar _gv_i_60;
											for (_gv_i_60 = 0; _gv_i_60 < BLOCK_SIZE; _gv_i_60 = _gv_i_60 + 1) begin : g_commit_in
												localparam i = _gv_i_60;
												// Trace: src/VX_gather_unit.sv:24:9
												assign result_in_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_result_if[i + _mbase_result_if].valid;
												// Trace: src/VX_gather_unit.sv:25:9
												assign result_in_data[i * 174+:174] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_result_if[i + _mbase_result_if].data;
												// Trace: src/VX_gather_unit.sv:26:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.alu_unit.per_block_result_if[i + _mbase_result_if].ready = result_in_ready[i];
												if (1) begin : g_result_in_isw_full
													// Trace: src/VX_gather_unit.sv:34:13
													assign result_in_isw[i+:1] = sv2v_cast_1_signed(i);
												end
											end
											// Trace: src/VX_gather_unit.sv:37:5
											reg [0:0] result_out_valid;
											// Trace: src/VX_gather_unit.sv:38:5
											reg [173:0] result_out_data;
											// Trace: src/VX_gather_unit.sv:39:5
											wire [0:0] result_out_ready;
											// Trace: src/VX_gather_unit.sv:40:5
											always @(*) begin
												// Trace: src/VX_gather_unit.sv:41:9
												result_out_valid = 1'sb0;
												// Trace: src/VX_gather_unit.sv:42:9
												begin : sv2v_autoblock_9
													// Trace: src/VX_gather_unit.sv:42:14
													integer i;
													// Trace: src/VX_gather_unit.sv:42:14
													for (i = 0; i < 1; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:43:13
															result_out_data[i * 174+:174] = 1'sbx;
														end
												end
												begin : sv2v_autoblock_10
													// Trace: src/VX_gather_unit.sv:45:14
													integer i;
													// Trace: src/VX_gather_unit.sv:45:14
													for (i = 0; i < BLOCK_SIZE; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:46:13
															result_out_valid[result_in_isw[i+:1]] = result_in_valid[i];
															// Trace: src/VX_gather_unit.sv:47:13
															result_out_data[result_in_isw[i+:1] * 174+:174] = result_in_data[i * 174+:174];
														end
												end
											end
											// Trace: src/VX_gather_unit.sv:50:5
											genvar _gv_i_61;
											for (_gv_i_61 = 0; _gv_i_61 < BLOCK_SIZE; _gv_i_61 = _gv_i_61 + 1) begin : g_result_in_ready
												localparam i = _gv_i_61;
												// Trace: src/VX_gather_unit.sv:51:9
												assign result_in_ready[i] = result_out_ready[result_in_isw[i+:1]];
											end
											// Trace: src/VX_gather_unit.sv:53:5
											genvar _gv_i_62;
											localparam VX_gpu_pkg_SIMD_COUNT = 1;
											localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
											localparam VX_gpu_pkg_SIMD_IDX_W = 1;
											for (_gv_i_62 = 0; _gv_i_62 < 1; _gv_i_62 = _gv_i_62 + 1) begin : g_out_bufs
												localparam i = _gv_i_62;
												// Trace: src/VX_gather_unit.sv:54:9
												// expanded interface instance: result_tmp_if
												localparam _param_D4A7C_NUM_LANES = NUM_LANES;
												if (1) begin : result_tmp_if
													// removed import VX_gpu_pkg::*;
													// Trace: src/VX_result_if.sv:2:15
													localparam NUM_LANES = _param_D4A7C_NUM_LANES;
													// Trace: src/VX_result_if.sv:3:15
													localparam PID_WIDTH = 1;
													// Trace: src/VX_result_if.sv:5:5
													localparam VX_gpu_pkg_REG_TYPES = 1;
													localparam VX_gpu_pkg_RV_REGS = 32;
													localparam VX_gpu_pkg_NUM_REGS = 32;
													localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
													localparam VX_gpu_pkg_NW_BITS = 2;
													localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
													localparam VX_gpu_pkg_PC_BITS = 30;
													localparam VX_gpu_pkg_UUID_WIDTH = 1;
													// removed localparam type data_t
													// Trace: src/VX_result_if.sv:17:5
													wire valid;
													// Trace: src/VX_result_if.sv:18:5
													wire [173:0] data;
													// Trace: src/VX_result_if.sv:19:5
													wire ready;
													// Trace: src/VX_result_if.sv:20:5
													// Trace: src/VX_result_if.sv:25:5
												end
												// Trace: src/VX_gather_unit.sv:57:9
												VX_elastic_buffer #(
													.DATAW(DATAW),
													.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
													.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
												) out_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(result_out_valid[i]),
													.ready_in(result_out_ready[i]),
													.data_in(result_out_data[i * 174+:174]),
													.data_out(result_tmp_if.data),
													.valid_out(result_tmp_if.valid),
													.ready_out(result_tmp_if.ready)
												);
												// Trace: src/VX_gather_unit.sv:71:9
												wire [0:0] commit_sid_w;
												// Trace: src/VX_gather_unit.sv:72:9
												wire [3:0] commit_tmask_w;
												// Trace: src/VX_gather_unit.sv:73:9
												wire [127:0] commit_data_w;
												if (1) begin : g_no_lpid
													// Trace: src/VX_gather_unit.sv:91:13
													assign commit_sid_w = result_tmp_if.data[2];
													// Trace: src/VX_gather_unit.sv:92:13
													assign commit_tmask_w = result_tmp_if.data[170-:4];
													// Trace: src/VX_gather_unit.sv:93:13
													assign commit_data_w = result_tmp_if.data[130-:128];
												end
												// Trace: src/VX_gather_unit.sv:95:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_if].valid = result_tmp_if.valid;
												// Trace: src/VX_gather_unit.sv:96:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_if].data = {result_tmp_if.data[173], result_tmp_if.data[172-:2], commit_sid_w, commit_tmask_w, result_tmp_if.data[166-:30], result_tmp_if.data[136], result_tmp_if.data[135-:5], commit_data_w, result_tmp_if.data[1], result_tmp_if.data[0]};
												// Trace: src/VX_gather_unit.sv:108:9
												assign result_tmp_if.ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_if].ready;
											end
										end
										assign gather_unit.clk = clk;
										assign gather_unit.reset = reset;
									end
									assign alu_unit.clk = clk;
									assign alu_unit.reset = reset;
									// Trace: src/VX_execute.sv:26:5
									localparam VX_gpu_pkg_EX_LSU = 1;
									// expanded module instance: lsu_unit
									localparam _bbase_54826_dispatch_if = 1;
									localparam _bbase_54826_commit_if = 1;
									localparam _bbase_54826_lsu_mem_if = 0;
									localparam _param_54826_INSTANCE_ID = "";
									if (1) begin : lsu_unit
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_lsu_unit.sv:2:15
										localparam INSTANCE_ID = _param_54826_INSTANCE_ID;
										// Trace: src/VX_lsu_unit.sv:4:5
										wire clk;
										// Trace: src/VX_lsu_unit.sv:5:5
										wire reset;
										// Trace: src/VX_lsu_unit.sv:6:5
										localparam _mbase_dispatch_if = 1;
										// Trace: src/VX_lsu_unit.sv:7:5
										localparam _mbase_commit_if = 1;
										// Trace: src/VX_lsu_unit.sv:8:5
										localparam _mbase_lsu_mem_if = 0;
										// Trace: src/VX_lsu_unit.sv:10:5
										localparam BLOCK_SIZE = 1;
										// Trace: src/VX_lsu_unit.sv:11:5
										localparam NUM_LANES = 4;
										// Trace: src/VX_lsu_unit.sv:13:5
										// expanded interface instance: per_block_execute_if
										localparam _param_E2592_NUM_LANES = NUM_LANES;
										genvar _arr_E2592;
										for (_arr_E2592 = 0; _arr_E2592 <= 0; _arr_E2592 = _arr_E2592 + 1) begin : per_block_execute_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_execute_if.sv:2:15
											localparam NUM_LANES = _param_E2592_NUM_LANES;
											// Trace: src/VX_execute_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_execute_if.sv:5:5
											localparam VX_gpu_pkg_INST_ALU_BITS = 4;
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
											// removed localparam type VX_gpu_pkg_alu_args_t
											localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
											// removed localparam type VX_gpu_pkg_csr_args_t
											localparam VX_gpu_pkg_INST_FMT_BITS = 2;
											localparam VX_gpu_pkg_INST_FRM_BITS = 3;
											// removed localparam type VX_gpu_pkg_fpu_args_t
											localparam VX_gpu_pkg_OFFSET_BITS = 12;
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											// removed localparam type data_t
											// Trace: src/VX_execute_if.sv:21:5
											wire valid;
											// Trace: src/VX_execute_if.sv:22:5
											wire [470:0] data;
											// Trace: src/VX_execute_if.sv:23:5
											wire ready;
											// Trace: src/VX_execute_if.sv:24:5
											// Trace: src/VX_execute_if.sv:29:5
										end
										// Trace: src/VX_lsu_unit.sv:16:5
										// expanded module instance: dispatch_unit
										localparam _bbase_2E16E_dispatch_if = 1;
										localparam _bbase_2E16E_execute_if = 0;
										localparam _param_2E16E_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_2E16E_NUM_LANES = NUM_LANES;
										localparam _param_2E16E_OUT_BUF = 3;
										if (1) begin : dispatch_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_dispatch_unit.sv:2:15
											localparam BLOCK_SIZE = _param_2E16E_BLOCK_SIZE;
											// Trace: src/VX_dispatch_unit.sv:3:15
											localparam NUM_LANES = _param_2E16E_NUM_LANES;
											// Trace: src/VX_dispatch_unit.sv:4:15
											localparam OUT_BUF = _param_2E16E_OUT_BUF;
											// Trace: src/VX_dispatch_unit.sv:5:15
											localparam MAX_FANOUT = 8;
											// Trace: src/VX_dispatch_unit.sv:7:5
											wire clk;
											// Trace: src/VX_dispatch_unit.sv:8:5
											wire reset;
											// Trace: src/VX_dispatch_unit.sv:9:5
											localparam _mbase_dispatch_if = 1;
											// Trace: src/VX_dispatch_unit.sv:10:5
											localparam _mbase_execute_if = 0;
											// Trace: src/VX_dispatch_unit.sv:12:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:13:5
											localparam NUM_PACKETS = 1;
											// Trace: src/VX_dispatch_unit.sv:14:5
											localparam LPID_BITS = 0;
											// Trace: src/VX_dispatch_unit.sv:15:5
											localparam LPID_WIDTH = 1;
											// Trace: src/VX_dispatch_unit.sv:16:5
											localparam GPID_BITS = 0;
											// Trace: src/VX_dispatch_unit.sv:17:5
											localparam GPID_WIDTH = 1;
											// Trace: src/VX_dispatch_unit.sv:18:5
											localparam BATCH_COUNT = 1;
											// Trace: src/VX_dispatch_unit.sv:19:5
											localparam BATCH_COUNT_W = 1;
											// Trace: src/VX_dispatch_unit.sv:20:5
											localparam ISSUE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:21:5
											localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
											localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
											localparam VX_gpu_pkg_INST_OP_BITS = 4;
											localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
											localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
											localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_SIMD_COUNT = 1;
											localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
											localparam VX_gpu_pkg_SIMD_IDX_W = 1;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam IN_DATAW = 471;
											// Trace: src/VX_dispatch_unit.sv:22:5
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam OUT_DATAW = 471;
											// Trace: src/VX_dispatch_unit.sv:23:5
											localparam FANOUT_ENABLE = 1'd0;
											// Trace: src/VX_dispatch_unit.sv:24:5
											localparam DATA_TMASK_OFF = 463;
											// Trace: src/VX_dispatch_unit.sv:25:5
											localparam DATA_REGS_OFF = 2;
											// Trace: src/VX_dispatch_unit.sv:26:5
											// removed localparam type packet_t
											// Trace: src/VX_dispatch_unit.sv:30:5
											wire [0:0] dispatch_valid;
											// Trace: src/VX_dispatch_unit.sv:31:5
											wire [470:0] dispatch_data;
											// Trace: src/VX_dispatch_unit.sv:32:5
											wire [0:0] dispatch_ready;
											// Trace: src/VX_dispatch_unit.sv:33:5
											genvar _gv_i_35;
											for (_gv_i_35 = 0; _gv_i_35 < 1; _gv_i_35 = _gv_i_35 + 1) begin : g_dispatch_data
												localparam i = _gv_i_35;
												// Trace: src/VX_dispatch_unit.sv:34:9
												assign dispatch_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].valid;
												// Trace: src/VX_dispatch_unit.sv:35:9
												assign dispatch_data[i * 471+:471] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].data;
												// Trace: src/VX_dispatch_unit.sv:36:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].ready = dispatch_ready[i];
											end
											// Trace: src/VX_dispatch_unit.sv:38:5
											wire [0:0] block_ready;
											// Trace: src/VX_dispatch_unit.sv:39:5
											wire [3:0] block_tmask;
											// Trace: src/VX_dispatch_unit.sv:40:5
											wire [383:0] block_rsdata;
											// Trace: src/VX_dispatch_unit.sv:41:5
											wire [0:0] block_pid;
											// Trace: src/VX_dispatch_unit.sv:42:5
											wire [0:0] block_sop;
											// Trace: src/VX_dispatch_unit.sv:43:5
											wire [0:0] block_eop;
											// Trace: src/VX_dispatch_unit.sv:44:5
											wire [0:0] block_done;
											// Trace: src/VX_dispatch_unit.sv:45:5
											wire batch_done = &block_done;
											// Trace: src/VX_dispatch_unit.sv:46:5
											wire [0:0] batch_idx;
											// Trace: src/VX_dispatch_unit.sv:47:5
											if (1) begin : g_batch_idx_0
												// Trace: src/VX_dispatch_unit.sv:73:9
												assign batch_idx = 0;
											end
											// Trace: src/VX_dispatch_unit.sv:75:5
											wire [0:0] issue_indices;
											// Trace: src/VX_dispatch_unit.sv:76:5
											genvar _gv_block_idx_2;
											for (_gv_block_idx_2 = 0; _gv_block_idx_2 < BLOCK_SIZE; _gv_block_idx_2 = _gv_block_idx_2 + 1) begin : g_issue_indices
												localparam block_idx = _gv_block_idx_2;
												// Trace: src/VX_dispatch_unit.sv:77:9
												assign issue_indices[block_idx+:1] = sv2v_cast_1(batch_idx * BLOCK_SIZE) + sv2v_cast_1_signed(block_idx);
											end
											// Trace: src/VX_dispatch_unit.sv:79:5
											genvar _gv_block_idx_3;
											localparam VX_gpu_pkg_ISSUE_ISW_BITS = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											function automatic [1:0] VX_gpu_pkg_wis_to_wid;
												// Trace: src/VX_gpu_pkg.sv:264:9
												input reg [1:0] wis;
												// Trace: src/VX_gpu_pkg.sv:265:9
												input reg [0:0] isw;
												// Trace: src/VX_gpu_pkg.sv:267:9
												begin
													// Trace: src/VX_gpu_pkg.sv:270:13
													VX_gpu_pkg_wis_to_wid = wis;
												end
											endfunction
											for (_gv_block_idx_3 = 0; _gv_block_idx_3 < BLOCK_SIZE; _gv_block_idx_3 = _gv_block_idx_3 + 1) begin : g_blocks
												localparam block_idx = _gv_block_idx_3;
												// Trace: src/VX_dispatch_unit.sv:80:9
												wire [0:0] issue_idx = issue_indices[block_idx+:1];
												// Trace: src/VX_dispatch_unit.sv:81:9
												wire [1:0] dispatch_wis = dispatch_data[(issue_idx * 471) + 468+:VX_gpu_pkg_ISSUE_WIS_W];
												// Trace: src/VX_dispatch_unit.sv:82:9
												wire [0:0] dispatch_sid = dispatch_data[(issue_idx * 471) + 467+:VX_gpu_pkg_SIMD_IDX_W];
												// Trace: src/VX_dispatch_unit.sv:83:9
												wire dispatch_sop = dispatch_data[(issue_idx * 471) + 1];
												// Trace: src/VX_dispatch_unit.sv:84:9
												wire dispatch_eop = dispatch_data[issue_idx * 471];
												// Trace: src/VX_dispatch_unit.sv:85:9
												wire [3:0] dispatch_tmask;
												// Trace: src/VX_dispatch_unit.sv:86:9
												wire [383:0] dispatch_rsdata;
												// Trace: src/VX_dispatch_unit.sv:87:9
												assign dispatch_tmask = dispatch_data[(issue_idx * 471) + DATA_TMASK_OFF+:4];
												// Trace: src/VX_dispatch_unit.sv:88:9
												assign dispatch_rsdata[0+:128] = dispatch_data[(issue_idx * 471) + 258+:128];
												// Trace: src/VX_dispatch_unit.sv:89:9
												assign dispatch_rsdata[128+:128] = dispatch_data[(issue_idx * 471) + 130+:128];
												// Trace: src/VX_dispatch_unit.sv:90:9
												assign dispatch_rsdata[256+:128] = dispatch_data[(issue_idx * 471) + 2+:128];
												// Trace: src/VX_dispatch_unit.sv:91:9
												wire valid_p;
												wire ready_p;
												if (1) begin : g_full_simd
													// Trace: src/VX_dispatch_unit.sv:132:13
													assign valid_p = dispatch_valid[issue_idx];
													// Trace: src/VX_dispatch_unit.sv:133:13
													assign block_tmask[block_idx * 4+:4] = dispatch_tmask;
													// Trace: src/VX_dispatch_unit.sv:134:13
													assign block_rsdata[32 * (4 * (block_idx * 3))+:384] = dispatch_rsdata;
													// Trace: src/VX_dispatch_unit.sv:135:13
													assign block_pid[block_idx+:1] = 0;
													// Trace: src/VX_dispatch_unit.sv:136:13
													assign block_sop[block_idx] = 1;
													// Trace: src/VX_dispatch_unit.sv:137:13
													assign block_eop[block_idx] = 1;
													// Trace: src/VX_dispatch_unit.sv:138:13
													assign block_ready[block_idx] = ready_p;
													// Trace: src/VX_dispatch_unit.sv:139:13
													assign block_done[block_idx] = ready_p || ~valid_p;
												end
												// Trace: src/VX_dispatch_unit.sv:141:9
												wire [0:0] isw;
												if (1) begin : g_isw
													// Trace: src/VX_dispatch_unit.sv:149:13
													assign isw = block_idx;
												end
												// Trace: src/VX_dispatch_unit.sv:151:9
												wire [1:0] block_wid = VX_gpu_pkg_wis_to_wid(dispatch_wis, isw);
												// Trace: src/VX_dispatch_unit.sv:152:9
												wire [0:0] warp_pid = block_pid[block_idx+:1] + sv2v_cast_1(dispatch_sid * NUM_PACKETS);
												// Trace: src/VX_dispatch_unit.sv:153:9
												wire warp_sop = block_sop[block_idx] && dispatch_sop;
												// Trace: src/VX_dispatch_unit.sv:154:9
												wire warp_eop = block_eop[block_idx] && dispatch_eop;
												// Trace: src/VX_dispatch_unit.sv:155:9
												VX_elastic_buffer #(
													.DATAW(OUT_DATAW),
													.SIZE(2),
													.OUT_REG(1)
												) buf_out(
													.clk(clk),
													.reset(reset),
													.valid_in(valid_p),
													.ready_in(ready_p),
													.data_in({dispatch_data[(issue_idx * 471) + 470-:VX_gpu_pkg_UUID_WIDTH], block_wid, block_tmask[block_idx * 4+:4], dispatch_data[(issue_idx * 471) + 462-:77], block_rsdata[32 * ((block_idx * 3) * 4)+:128], block_rsdata[32 * (((block_idx * 3) + 1) * 4)+:128], block_rsdata[32 * (((block_idx * 3) + 2) * 4)+:128], warp_pid, warp_sop, warp_eop}),
													.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[block_idx + _mbase_execute_if].data),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[block_idx + _mbase_execute_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[block_idx + _mbase_execute_if].ready)
												);
											end
											// Trace: src/VX_dispatch_unit.sv:180:5
											reg [0:0] ready_in;
											// Trace: src/VX_dispatch_unit.sv:181:5
											always @(*) begin
												// Trace: src/VX_dispatch_unit.sv:182:9
												ready_in = 0;
												// Trace: src/VX_dispatch_unit.sv:183:9
												begin : sv2v_autoblock_11
													// Trace: src/VX_dispatch_unit.sv:183:14
													integer block_idx;
													// Trace: src/VX_dispatch_unit.sv:183:14
													for (block_idx = 0; block_idx < BLOCK_SIZE; block_idx = block_idx + 1)
														begin
															// Trace: src/VX_dispatch_unit.sv:184:13
															ready_in[issue_indices[block_idx+:1]] = block_ready[block_idx] && block_eop[block_idx];
														end
												end
											end
											// Trace: src/VX_dispatch_unit.sv:187:5
											assign dispatch_ready = ready_in;
										end
										assign dispatch_unit.clk = clk;
										assign dispatch_unit.reset = reset;
										// Trace: src/VX_lsu_unit.sv:26:5
										// expanded interface instance: per_block_result_if
										localparam _param_911F6_NUM_LANES = NUM_LANES;
										genvar _arr_911F6;
										for (_arr_911F6 = 0; _arr_911F6 <= 0; _arr_911F6 = _arr_911F6 + 1) begin : per_block_result_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_result_if.sv:2:15
											localparam NUM_LANES = _param_911F6_NUM_LANES;
											// Trace: src/VX_result_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_result_if.sv:5:5
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											// removed localparam type data_t
											// Trace: src/VX_result_if.sv:17:5
											wire valid;
											// Trace: src/VX_result_if.sv:18:5
											wire [173:0] data;
											// Trace: src/VX_result_if.sv:19:5
											wire ready;
											// Trace: src/VX_result_if.sv:20:5
											// Trace: src/VX_result_if.sv:25:5
										end
										// Trace: src/VX_lsu_unit.sv:29:5
										genvar _gv_block_idx_5;
										for (_gv_block_idx_5 = 0; _gv_block_idx_5 < BLOCK_SIZE; _gv_block_idx_5 = _gv_block_idx_5 + 1) begin : g_blocks
											localparam block_idx = _gv_block_idx_5;
											// Trace: src/VX_lsu_unit.sv:30:9
											// expanded module instance: lsu_slice
											localparam _bbase_DE6D2_execute_if = block_idx;
											localparam _bbase_DE6D2_result_if = block_idx;
											localparam _bbase_DE6D2_lsu_mem_if = block_idx + _mbase_lsu_mem_if;
											localparam _param_DE6D2_INSTANCE_ID = "";
											if (1) begin : lsu_slice
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_lsu_slice.sv:2:15
												localparam INSTANCE_ID = _param_DE6D2_INSTANCE_ID;
												// Trace: src/VX_lsu_slice.sv:4:5
												wire clk;
												// Trace: src/VX_lsu_slice.sv:5:5
												wire reset;
												// Trace: src/VX_lsu_slice.sv:6:5
												localparam _mbase_execute_if = _bbase_DE6D2_execute_if;
												// Trace: src/VX_lsu_slice.sv:7:5
												localparam _mbase_result_if = _bbase_DE6D2_result_if;
												// Trace: src/VX_lsu_slice.sv:8:5
												localparam _mbase_lsu_mem_if = _bbase_DE6D2_lsu_mem_if;
												// Trace: src/VX_lsu_slice.sv:10:5
												localparam NUM_LANES = 4;
												// Trace: src/VX_lsu_slice.sv:11:5
												localparam PID_BITS = 0;
												// Trace: src/VX_lsu_slice.sv:12:5
												localparam PID_WIDTH = 1;
												// Trace: src/VX_lsu_slice.sv:13:5
												localparam VX_gpu_pkg_REG_TYPES = 1;
												localparam VX_gpu_pkg_RV_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS = 32;
												localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
												localparam VX_gpu_pkg_NW_BITS = 2;
												localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
												localparam VX_gpu_pkg_PC_BITS = 30;
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												localparam RSP_ARB_DATAW = 174;
												// Trace: src/VX_lsu_slice.sv:14:5
												localparam LSUQ_SIZEW = 1;
												// Trace: src/VX_lsu_slice.sv:15:5
												localparam VX_gpu_pkg_XLENB = 4;
												localparam VX_gpu_pkg_LSU_WORD_SIZE = VX_gpu_pkg_XLENB;
												localparam REQ_ASHIFT = 2;
												// Trace: src/VX_lsu_slice.sv:16:5
												localparam MEM_ASHIFT = 6;
												// Trace: src/VX_lsu_slice.sv:17:5
												localparam MEM_ADDRW = 26;
												// Trace: src/VX_lsu_slice.sv:18:5
												localparam VX_gpu_pkg_INST_LSU_BITS = 4;
												localparam TAG_ID_WIDTH = 53;
												// Trace: src/VX_lsu_slice.sv:19:5
												localparam TAG_WIDTH = 54;
												// Trace: src/VX_lsu_slice.sv:20:5
												// expanded interface instance: result_rsp_if
												localparam _param_3E3A8_NUM_LANES = NUM_LANES;
												if (1) begin : result_rsp_if
													// removed import VX_gpu_pkg::*;
													// Trace: src/VX_result_if.sv:2:15
													localparam NUM_LANES = _param_3E3A8_NUM_LANES;
													// Trace: src/VX_result_if.sv:3:15
													localparam PID_WIDTH = 1;
													// Trace: src/VX_result_if.sv:5:5
													localparam VX_gpu_pkg_REG_TYPES = 1;
													localparam VX_gpu_pkg_RV_REGS = 32;
													localparam VX_gpu_pkg_NUM_REGS = 32;
													localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
													localparam VX_gpu_pkg_NW_BITS = 2;
													localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
													localparam VX_gpu_pkg_PC_BITS = 30;
													localparam VX_gpu_pkg_UUID_WIDTH = 1;
													// removed localparam type data_t
													// Trace: src/VX_result_if.sv:17:5
													wire valid;
													// Trace: src/VX_result_if.sv:18:5
													wire [173:0] data;
													// Trace: src/VX_result_if.sv:19:5
													wire ready;
													// Trace: src/VX_result_if.sv:20:5
													// Trace: src/VX_result_if.sv:25:5
												end
												// Trace: src/VX_lsu_slice.sv:23:5
												// expanded interface instance: result_no_rsp_if
												localparam _param_B28AB_NUM_LANES = NUM_LANES;
												if (1) begin : result_no_rsp_if
													// removed import VX_gpu_pkg::*;
													// Trace: src/VX_result_if.sv:2:15
													localparam NUM_LANES = _param_B28AB_NUM_LANES;
													// Trace: src/VX_result_if.sv:3:15
													localparam PID_WIDTH = 1;
													// Trace: src/VX_result_if.sv:5:5
													localparam VX_gpu_pkg_REG_TYPES = 1;
													localparam VX_gpu_pkg_RV_REGS = 32;
													localparam VX_gpu_pkg_NUM_REGS = 32;
													localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
													localparam VX_gpu_pkg_NW_BITS = 2;
													localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
													localparam VX_gpu_pkg_PC_BITS = 30;
													localparam VX_gpu_pkg_UUID_WIDTH = 1;
													// removed localparam type data_t
													// Trace: src/VX_result_if.sv:17:5
													wire valid;
													// Trace: src/VX_result_if.sv:18:5
													wire [173:0] data;
													// Trace: src/VX_result_if.sv:19:5
													wire ready;
													// Trace: src/VX_result_if.sv:20:5
													// Trace: src/VX_result_if.sv:25:5
												end
												// Trace: src/VX_lsu_slice.sv:26:5
												wire req_is_fence;
												wire rsp_is_fence;
												// Trace: src/VX_lsu_slice.sv:27:5
												wire [127:0] full_addr;
												// Trace: src/VX_lsu_slice.sv:28:5
												genvar _gv_i_113;
												for (_gv_i_113 = 0; _gv_i_113 < NUM_LANES; _gv_i_113 = _gv_i_113 + 1) begin : g_full_addr
													localparam i = _gv_i_113;
													// Trace: src/VX_lsu_slice.sv:29:9
													assign full_addr[i * 32+:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[259 + (i * 32)+:32] + {{21 {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[404]}}, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[403:393]};
												end
												// Trace: src/VX_lsu_slice.sv:31:5
												localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
												localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
												wire [11:0] mem_req_flags;
												// Trace: src/VX_lsu_slice.sv:32:5
												genvar _gv_i_114;
												localparam VX_gpu_pkg_MEM_REQ_FLAG_FLUSH = 0;
												localparam VX_gpu_pkg_MEM_REQ_FLAG_IO = 1;
												for (_gv_i_114 = 0; _gv_i_114 < NUM_LANES; _gv_i_114 = _gv_i_114 + 1) begin : g_mem_req_flags
													localparam i = _gv_i_114;
													// Trace: src/VX_lsu_slice.sv:33:9
													wire [25:0] block_addr = full_addr[(i * 32) + MEM_ASHIFT+:MEM_ADDRW];
													// Trace: src/VX_lsu_slice.sv:34:9
													wire [25:0] io_addr_start = sv2v_cast_26(32'h00000040 >> MEM_ASHIFT);
													// Trace: src/VX_lsu_slice.sv:35:9
													wire [25:0] io_addr_end = sv2v_cast_26(32'h00010000 >> MEM_ASHIFT);
													// Trace: src/VX_lsu_slice.sv:36:9
													assign mem_req_flags[(i * 3) + VX_gpu_pkg_MEM_REQ_FLAG_FLUSH] = req_is_fence;
													// Trace: src/VX_lsu_slice.sv:37:9
													assign mem_req_flags[(i * 3) + VX_gpu_pkg_MEM_REQ_FLAG_IO] = (block_addr >= io_addr_start) && (block_addr < io_addr_end);
													// Trace: src/VX_lsu_slice.sv:38:9
													wire [25:0] lmem_addr_start = sv2v_cast_26(32'hffff0000 >> MEM_ASHIFT);
													// Trace: src/VX_lsu_slice.sv:39:9
													wire [25:0] lmem_addr_end = sv2v_cast_26((32'hffff0000 + 32'sd16384) >> MEM_ASHIFT);
													// Trace: src/VX_lsu_slice.sv:40:9
													assign mem_req_flags[(i * 3) + VX_gpu_pkg_MEM_REQ_FLAG_LOCAL] = (block_addr >= lmem_addr_start) && (block_addr < lmem_addr_end);
												end
												// Trace: src/VX_lsu_slice.sv:42:5
												wire mem_req_valid;
												// Trace: src/VX_lsu_slice.sv:43:5
												wire [3:0] mem_req_mask;
												// Trace: src/VX_lsu_slice.sv:44:5
												wire mem_req_rw;
												// Trace: src/VX_lsu_slice.sv:45:5
												localparam VX_gpu_pkg_LSU_ADDR_WIDTH = 30;
												wire [119:0] mem_req_addr;
												// Trace: src/VX_lsu_slice.sv:46:5
												wire [15:0] mem_req_byteen;
												// Trace: src/VX_lsu_slice.sv:47:5
												reg [127:0] mem_req_data;
												// Trace: src/VX_lsu_slice.sv:48:5
												wire [53:0] mem_req_tag;
												// Trace: src/VX_lsu_slice.sv:49:5
												wire mem_req_ready;
												// Trace: src/VX_lsu_slice.sv:50:5
												wire mem_rsp_valid;
												// Trace: src/VX_lsu_slice.sv:51:5
												wire [3:0] mem_rsp_mask;
												// Trace: src/VX_lsu_slice.sv:52:5
												wire [127:0] mem_rsp_data;
												// Trace: src/VX_lsu_slice.sv:53:5
												wire [53:0] mem_rsp_tag;
												// Trace: src/VX_lsu_slice.sv:54:5
												wire mem_rsp_sop;
												// Trace: src/VX_lsu_slice.sv:55:5
												wire mem_rsp_eop;
												// Trace: src/VX_lsu_slice.sv:56:5
												wire mem_rsp_ready;
												// Trace: src/VX_lsu_slice.sv:57:5
												wire mem_req_fire = mem_req_valid && mem_req_ready;
												// Trace: src/VX_lsu_slice.sv:58:5
												wire mem_rsp_fire = mem_rsp_valid && mem_rsp_ready;
												// Trace: src/VX_lsu_slice.sv:59:5
												wire mem_rsp_sop_pkt;
												wire mem_rsp_eop_pkt;
												// Trace: src/VX_lsu_slice.sv:60:5
												wire no_rsp_buf_valid;
												wire no_rsp_buf_ready;
												// Trace: src/VX_lsu_slice.sv:61:5
												wire [0:0] pkt_waddr;
												wire [0:0] pkt_raddr;
												// Trace: src/VX_lsu_slice.sv:62:5
												reg fence_lock;
												// Trace: src/VX_lsu_slice.sv:63:5
												function automatic VX_gpu_pkg_inst_lsu_is_fence;
													// Trace: src/VX_gpu_pkg.sv:216:48
													input reg [3:0] op;
													// Trace: src/VX_gpu_pkg.sv:217:9
													VX_gpu_pkg_inst_lsu_is_fence = op[3:2] == 3;
												endfunction
												assign req_is_fence = VX_gpu_pkg_inst_lsu_is_fence(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[433-:4]);
												// Trace: src/VX_lsu_slice.sv:64:5
												always @(posedge clk)
													// Trace: src/VX_lsu_slice.sv:65:9
													if (reset)
														// Trace: src/VX_lsu_slice.sv:66:13
														fence_lock <= 0;
													else begin
														// Trace: src/VX_lsu_slice.sv:68:13
														if ((mem_req_fire && req_is_fence) && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[0])
															// Trace: src/VX_lsu_slice.sv:69:17
															fence_lock <= 1;
														if ((mem_rsp_fire && rsp_is_fence) && mem_rsp_eop_pkt)
															// Trace: src/VX_lsu_slice.sv:72:17
															fence_lock <= 0;
													end
												// Trace: src/VX_lsu_slice.sv:76:5
												wire req_skip = req_is_fence && ~Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[0];
												// Trace: src/VX_lsu_slice.sv:77:5
												wire no_rsp_buf_enable = (mem_req_rw && ~Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[392]) || req_skip;
												// Trace: src/VX_lsu_slice.sv:78:5
												assign mem_req_valid = ((Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].valid && ~req_skip) && ~(no_rsp_buf_enable && ~no_rsp_buf_ready)) && ~fence_lock;
												// Trace: src/VX_lsu_slice.sv:82:5
												assign no_rsp_buf_valid = ((Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].valid && no_rsp_buf_enable) && (req_skip || mem_req_ready)) && ~fence_lock;
												// Trace: src/VX_lsu_slice.sv:86:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].ready = ((mem_req_ready || req_skip) && ~(no_rsp_buf_enable && ~no_rsp_buf_ready)) && ~fence_lock;
												// Trace: src/VX_lsu_slice.sv:89:5
												assign mem_req_mask = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[467-:4];
												// Trace: src/VX_lsu_slice.sv:90:5
												assign mem_req_rw = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[406];
												// Trace: src/VX_lsu_slice.sv:91:5
												wire [7:0] req_align;
												// Trace: src/VX_lsu_slice.sv:92:5
												genvar _gv_i_115;
												for (_gv_i_115 = 0; _gv_i_115 < NUM_LANES; _gv_i_115 = _gv_i_115 + 1) begin : g_mem_req_addr
													localparam i = _gv_i_115;
													// Trace: src/VX_lsu_slice.sv:93:9
													assign req_align[i * 2+:2] = full_addr[(i * 32) + 1-:2];
													// Trace: src/VX_lsu_slice.sv:94:9
													assign mem_req_addr[i * 30+:30] = full_addr[(i * 32) + 31-:30];
												end
												// Trace: src/VX_lsu_slice.sv:96:5
												genvar _gv_i_116;
												function automatic [1:0] VX_gpu_pkg_inst_lsu_wsize;
													// Trace: src/VX_gpu_pkg.sv:213:51
													input reg [3:0] op;
													// Trace: src/VX_gpu_pkg.sv:214:9
													VX_gpu_pkg_inst_lsu_wsize = op[1:0];
												endfunction
												for (_gv_i_116 = 0; _gv_i_116 < NUM_LANES; _gv_i_116 = _gv_i_116 + 1) begin : g_mem_req_byteen_w
													localparam i = _gv_i_116;
													// Trace: src/VX_lsu_slice.sv:97:9
													reg [3:0] mem_req_byteen_w;
													// Trace: src/VX_lsu_slice.sv:98:9
													always @(*) begin
														// Trace: src/VX_lsu_slice.sv:99:13
														mem_req_byteen_w = 1'sb0;
														// Trace: src/VX_lsu_slice.sv:100:13
														case (VX_gpu_pkg_inst_lsu_wsize(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[433-:4]))
															0:
																// Trace: src/VX_lsu_slice.sv:102:21
																mem_req_byteen_w[req_align[i * 2+:2]] = 1'b1;
															1: begin
																// Trace: src/VX_lsu_slice.sv:105:21
																mem_req_byteen_w[{req_align[(i * 2) + 1-:1], 1'b0}] = 1'b1;
																// Trace: src/VX_lsu_slice.sv:106:21
																mem_req_byteen_w[{req_align[(i * 2) + 1-:1], 1'b1}] = 1'b1;
															end
															default:
																// Trace: src/VX_lsu_slice.sv:108:27
																mem_req_byteen_w = {VX_gpu_pkg_LSU_WORD_SIZE {1'b1}};
														endcase
													end
													// Trace: src/VX_lsu_slice.sv:111:9
													assign mem_req_byteen[i * 4+:4] = mem_req_byteen_w;
												end
												// Trace: src/VX_lsu_slice.sv:113:5
												genvar _gv_i_117;
												for (_gv_i_117 = 0; _gv_i_117 < NUM_LANES; _gv_i_117 = _gv_i_117 + 1) begin : g_missalign
													localparam i = _gv_i_117;
													// Trace: src/VX_lsu_slice.sv:114:9
													wire lsu_req_fire = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].ready;
												end
												// Trace: src/VX_lsu_slice.sv:116:5
												genvar _gv_i_118;
												for (_gv_i_118 = 0; _gv_i_118 < NUM_LANES; _gv_i_118 = _gv_i_118 + 1) begin : g_mem_req_data
													localparam i = _gv_i_118;
													// Trace: src/VX_lsu_slice.sv:117:9
													always @(*) begin
														// Trace: src/VX_lsu_slice.sv:118:13
														mem_req_data[i * 32+:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[131 + (i * 32)+:32];
														// Trace: src/VX_lsu_slice.sv:119:13
														case (req_align[i * 2+:2])
															1:
																// Trace: src/VX_lsu_slice.sv:120:20
																mem_req_data[(i * 32) + 31-:24] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[131 + ((i * 32) + 23)-:24];
															2:
																// Trace: src/VX_lsu_slice.sv:121:20
																mem_req_data[(i * 32) + 31-:16] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[131 + ((i * 32) + 15)-:16];
															3:
																// Trace: src/VX_lsu_slice.sv:122:20
																mem_req_data[(i * 32) + 31-:8] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[131 + ((i * 32) + 7)-:8];
															default:
																;
														endcase
													end
												end
												// Trace: src/VX_lsu_slice.sv:127:5
												if (1) begin : g_no_pid
													// Trace: src/VX_lsu_slice.sv:180:9
													assign pkt_waddr = 0;
													// Trace: src/VX_lsu_slice.sv:181:9
													assign mem_rsp_sop_pkt = mem_rsp_sop;
													// Trace: src/VX_lsu_slice.sv:182:9
													assign mem_rsp_eop_pkt = mem_rsp_eop;
												end
												// Trace: src/VX_lsu_slice.sv:184:5
												assign mem_req_tag = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[470], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[469-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[463-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[392], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[391-:5], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[433-:4], req_align, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[2], pkt_waddr, req_is_fence};
												// Trace: src/VX_lsu_slice.sv:196:5
												wire lsu_mem_req_valid;
												// Trace: src/VX_lsu_slice.sv:197:5
												wire lsu_mem_req_rw;
												// Trace: src/VX_lsu_slice.sv:198:5
												wire [3:0] lsu_mem_req_mask;
												// Trace: src/VX_lsu_slice.sv:199:5
												wire [15:0] lsu_mem_req_byteen;
												// Trace: src/VX_lsu_slice.sv:200:5
												wire [119:0] lsu_mem_req_addr;
												// Trace: src/VX_lsu_slice.sv:201:5
												wire [11:0] lsu_mem_req_flags;
												// Trace: src/VX_lsu_slice.sv:202:5
												wire [127:0] lsu_mem_req_data;
												// Trace: src/VX_lsu_slice.sv:203:5
												localparam VX_gpu_pkg_LSU_MEM_BATCHES = 1;
												localparam VX_gpu_pkg_LSU_TAG_ID_BITS = 1;
												localparam VX_gpu_pkg_LSU_TAG_WIDTH = 2;
												wire [1:0] lsu_mem_req_tag;
												// Trace: src/VX_lsu_slice.sv:204:5
												wire lsu_mem_req_ready;
												// Trace: src/VX_lsu_slice.sv:205:5
												wire lsu_mem_rsp_valid;
												// Trace: src/VX_lsu_slice.sv:206:5
												wire [3:0] lsu_mem_rsp_mask;
												// Trace: src/VX_lsu_slice.sv:207:5
												wire [127:0] lsu_mem_rsp_data;
												// Trace: src/VX_lsu_slice.sv:208:5
												wire [1:0] lsu_mem_rsp_tag;
												// Trace: src/VX_lsu_slice.sv:209:5
												wire lsu_mem_rsp_ready;
												// Trace: src/VX_lsu_slice.sv:210:5
												VX_mem_scheduler #(
													.INSTANCE_ID(""),
													.CORE_REQS(NUM_LANES),
													.MEM_CHANNELS(NUM_LANES),
													.WORD_SIZE(VX_gpu_pkg_LSU_WORD_SIZE),
													.LINE_SIZE(VX_gpu_pkg_LSU_WORD_SIZE),
													.ADDR_WIDTH(VX_gpu_pkg_LSU_ADDR_WIDTH),
													.FLAGS_WIDTH(VX_gpu_pkg_MEM_FLAGS_WIDTH),
													.TAG_WIDTH(TAG_WIDTH),
													.CORE_QUEUE_SIZE(2),
													.MEM_QUEUE_SIZE(4),
													.UUID_WIDTH(VX_gpu_pkg_UUID_WIDTH),
													.RSP_PARTIAL(1),
													.MEM_OUT_BUF(0),
													.CORE_OUT_BUF(0)
												) mem_scheduler(
													.clk(clk),
													.reset(reset),
													.core_req_valid(mem_req_valid),
													.core_req_rw(mem_req_rw),
													.core_req_mask(mem_req_mask),
													.core_req_byteen(mem_req_byteen),
													.core_req_addr(mem_req_addr),
													.core_req_flags(mem_req_flags),
													.core_req_data(mem_req_data),
													.core_req_tag(mem_req_tag),
													.core_req_ready(mem_req_ready),
													.req_queue_empty(),
													.req_queue_rw_notify(),
													.core_rsp_valid(mem_rsp_valid),
													.core_rsp_mask(mem_rsp_mask),
													.core_rsp_data(mem_rsp_data),
													.core_rsp_tag(mem_rsp_tag),
													.core_rsp_sop(mem_rsp_sop),
													.core_rsp_eop(mem_rsp_eop),
													.core_rsp_ready(mem_rsp_ready),
													.mem_req_valid(lsu_mem_req_valid),
													.mem_req_rw(lsu_mem_req_rw),
													.mem_req_mask(lsu_mem_req_mask),
													.mem_req_byteen(lsu_mem_req_byteen),
													.mem_req_addr(lsu_mem_req_addr),
													.mem_req_flags(lsu_mem_req_flags),
													.mem_req_data(lsu_mem_req_data),
													.mem_req_tag(lsu_mem_req_tag),
													.mem_req_ready(lsu_mem_req_ready),
													.mem_rsp_valid(lsu_mem_rsp_valid),
													.mem_rsp_mask(lsu_mem_rsp_mask),
													.mem_rsp_data(lsu_mem_rsp_data),
													.mem_rsp_tag(lsu_mem_rsp_tag),
													.mem_rsp_ready(lsu_mem_rsp_ready)
												);
												// Trace: src/VX_lsu_slice.sv:261:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_valid = lsu_mem_req_valid;
												// Trace: src/VX_lsu_slice.sv:262:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[282-:4] = lsu_mem_req_mask;
												// Trace: src/VX_lsu_slice.sv:263:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[278] = lsu_mem_req_rw;
												// Trace: src/VX_lsu_slice.sv:264:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[29-:16] = lsu_mem_req_byteen;
												// Trace: src/VX_lsu_slice.sv:265:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[277-:120] = lsu_mem_req_addr;
												// Trace: src/VX_lsu_slice.sv:266:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[13-:12] = lsu_mem_req_flags;
												// Trace: src/VX_lsu_slice.sv:267:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[157-:128] = lsu_mem_req_data;
												// Trace: src/VX_lsu_slice.sv:268:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_data[1-:2] = lsu_mem_req_tag;
												// Trace: src/VX_lsu_slice.sv:269:5
												assign lsu_mem_req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].req_ready;
												// Trace: src/VX_lsu_slice.sv:270:5
												assign lsu_mem_rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].rsp_valid;
												// Trace: src/VX_lsu_slice.sv:271:5
												assign lsu_mem_rsp_mask = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].rsp_data[133-:4];
												// Trace: src/VX_lsu_slice.sv:272:5
												assign lsu_mem_rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].rsp_data[129-:128];
												// Trace: src/VX_lsu_slice.sv:273:5
												assign lsu_mem_rsp_tag = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].rsp_data[1-:2];
												// Trace: src/VX_lsu_slice.sv:274:5
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_mem_if].rsp_ready = lsu_mem_rsp_ready;
												// Trace: src/VX_lsu_slice.sv:275:5
												wire [0:0] rsp_uuid;
												// Trace: src/VX_lsu_slice.sv:276:5
												wire [1:0] rsp_wid;
												// Trace: src/VX_lsu_slice.sv:277:5
												wire [29:0] rsp_pc;
												// Trace: src/VX_lsu_slice.sv:278:5
												wire rsp_wb;
												// Trace: src/VX_lsu_slice.sv:279:5
												wire [4:0] rsp_rd;
												// Trace: src/VX_lsu_slice.sv:280:5
												wire [3:0] rsp_op_type;
												// Trace: src/VX_lsu_slice.sv:281:5
												wire [7:0] rsp_align;
												// Trace: src/VX_lsu_slice.sv:282:5
												wire [0:0] rsp_pid;
												// Trace: src/VX_lsu_slice.sv:283:5
												assign {rsp_uuid, rsp_wid, rsp_pc, rsp_wb, rsp_rd, rsp_op_type, rsp_align, rsp_pid, pkt_raddr, rsp_is_fence} = mem_rsp_tag;
												// Trace: src/VX_lsu_slice.sv:295:5
												reg [127:0] rsp_data;
												// Trace: src/VX_lsu_slice.sv:296:5
												genvar _gv_i_119;
												localparam VX_gpu_pkg_LSU_FMT_B = 3'b000;
												localparam VX_gpu_pkg_LSU_FMT_BU = 3'b100;
												localparam VX_gpu_pkg_LSU_FMT_H = 3'b001;
												localparam VX_gpu_pkg_LSU_FMT_HU = 3'b101;
												localparam VX_gpu_pkg_LSU_FMT_W = 3'b010;
												function automatic [2:0] VX_gpu_pkg_inst_lsu_fmt;
													// Trace: src/VX_gpu_pkg.sv:210:49
													input reg [3:0] op;
													// Trace: src/VX_gpu_pkg.sv:211:9
													VX_gpu_pkg_inst_lsu_fmt = op[2:0];
												endfunction
												for (_gv_i_119 = 0; _gv_i_119 < NUM_LANES; _gv_i_119 = _gv_i_119 + 1) begin : g_rsp_data
													localparam i = _gv_i_119;
													// Trace: src/VX_lsu_slice.sv:297:9
													wire [31:0] rsp_data32 = mem_rsp_data[i * 32+:32];
													// Trace: src/VX_lsu_slice.sv:298:9
													wire [15:0] rsp_data16 = (rsp_align[(i * 2) + 1] ? rsp_data32[31:16] : rsp_data32[15:0]);
													// Trace: src/VX_lsu_slice.sv:299:9
													wire [7:0] rsp_data8 = (rsp_align[i * 2] ? rsp_data16[15:8] : rsp_data16[7:0]);
													// Trace: src/VX_lsu_slice.sv:300:9
													always @(*)
														// Trace: src/VX_lsu_slice.sv:301:13
														case (VX_gpu_pkg_inst_lsu_fmt(rsp_op_type))
															VX_gpu_pkg_LSU_FMT_B:
																// Trace: src/VX_lsu_slice.sv:302:25
																rsp_data[i * 32+:32] = sv2v_cast_32_signed($signed(rsp_data8));
															VX_gpu_pkg_LSU_FMT_H:
																// Trace: src/VX_lsu_slice.sv:303:25
																rsp_data[i * 32+:32] = sv2v_cast_32_signed($signed(rsp_data16));
															VX_gpu_pkg_LSU_FMT_BU:
																// Trace: src/VX_lsu_slice.sv:304:25
																rsp_data[i * 32+:32] = sv2v_cast_32($unsigned(rsp_data8));
															VX_gpu_pkg_LSU_FMT_HU:
																// Trace: src/VX_lsu_slice.sv:305:25
																rsp_data[i * 32+:32] = sv2v_cast_32($unsigned(rsp_data16));
															VX_gpu_pkg_LSU_FMT_W:
																// Trace: src/VX_lsu_slice.sv:306:25
																rsp_data[i * 32+:32] = sv2v_cast_32_signed($signed(rsp_data32));
															default:
																// Trace: src/VX_lsu_slice.sv:307:22
																rsp_data[i * 32+:32] = 1'sbx;
														endcase
												end
												// Trace: src/VX_lsu_slice.sv:311:5
												VX_elastic_buffer #(
													.DATAW(174),
													.SIZE(2)
												) rsp_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(mem_rsp_valid),
													.ready_in(mem_rsp_ready),
													.data_in({rsp_uuid, rsp_wid, mem_rsp_mask, rsp_pc, rsp_wb, rsp_rd, rsp_data, rsp_pid, mem_rsp_sop_pkt, mem_rsp_eop_pkt}),
													.data_out({result_rsp_if.data[173], result_rsp_if.data[172-:2], result_rsp_if.data[170-:4], result_rsp_if.data[166-:30], result_rsp_if.data[136], result_rsp_if.data[135-:5], result_rsp_if.data[130-:128], result_rsp_if.data[2], result_rsp_if.data[1], result_rsp_if.data[0]}),
													.valid_out(result_rsp_if.valid),
													.ready_out(result_rsp_if.ready)
												);
												// Trace: src/VX_lsu_slice.sv:324:5
												VX_elastic_buffer #(
													.DATAW(40),
													.SIZE(2)
												) no_rsp_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(no_rsp_buf_valid),
													.ready_in(no_rsp_buf_ready),
													.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[470], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[469-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[467-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[463-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_execute_if[_mbase_execute_if].data[0]}),
													.data_out({result_no_rsp_if.data[173], result_no_rsp_if.data[172-:2], result_no_rsp_if.data[170-:4], result_no_rsp_if.data[166-:30], result_no_rsp_if.data[2], result_no_rsp_if.data[1], result_no_rsp_if.data[0]}),
													.valid_out(result_no_rsp_if.valid),
													.ready_out(result_no_rsp_if.ready)
												);
												// Trace: src/VX_lsu_slice.sv:337:5
												assign result_no_rsp_if.data[135-:5] = 1'sb0;
												// Trace: src/VX_lsu_slice.sv:338:5
												assign result_no_rsp_if.data[136] = 1'b0;
												// Trace: src/VX_lsu_slice.sv:339:5
												assign result_no_rsp_if.data[130-:128] = result_rsp_if.data[130-:128];
												// Trace: src/VX_lsu_slice.sv:340:5
												VX_stream_arb #(
													.NUM_INPUTS(2),
													.DATAW(RSP_ARB_DATAW),
													.ARBITER("P"),
													.OUT_BUF(3)
												) rsp_arb(
													.clk(clk),
													.reset(reset),
													.valid_in({result_no_rsp_if.valid, result_rsp_if.valid}),
													.ready_in({result_no_rsp_if.ready, result_rsp_if.ready}),
													.data_in({result_no_rsp_if.data, result_rsp_if.data}),
													.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_result_if[_mbase_result_if].data),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_result_if[_mbase_result_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_result_if[_mbase_result_if].ready),
													.sel_out()
												);
											end
											assign lsu_slice.clk = clk;
											assign lsu_slice.reset = reset;
										end
										// Trace: src/VX_lsu_unit.sv:40:5
										// expanded module instance: gather_unit
										localparam _bbase_8E516_result_if = 0;
										localparam _bbase_8E516_commit_if = 1;
										localparam _param_8E516_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_8E516_NUM_LANES = NUM_LANES;
										localparam _param_8E516_OUT_BUF = 3;
										if (1) begin : gather_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_gather_unit.sv:2:15
											localparam BLOCK_SIZE = _param_8E516_BLOCK_SIZE;
											// Trace: src/VX_gather_unit.sv:3:15
											localparam NUM_LANES = _param_8E516_NUM_LANES;
											// Trace: src/VX_gather_unit.sv:4:15
											localparam OUT_BUF = _param_8E516_OUT_BUF;
											// Trace: src/VX_gather_unit.sv:6:5
											wire clk;
											// Trace: src/VX_gather_unit.sv:7:5
											wire reset;
											// Trace: src/VX_gather_unit.sv:8:5
											localparam _mbase_result_if = 0;
											// Trace: src/VX_gather_unit.sv:9:5
											localparam _mbase_commit_if = 1;
											// Trace: src/VX_gather_unit.sv:11:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_gather_unit.sv:12:5
											localparam NUM_PACKETS = 1;
											// Trace: src/VX_gather_unit.sv:13:5
											localparam LPID_BITS = 0;
											// Trace: src/VX_gather_unit.sv:14:5
											localparam LPID_WIDTH = 1;
											// Trace: src/VX_gather_unit.sv:15:5
											localparam GPID_BITS = 0;
											// Trace: src/VX_gather_unit.sv:16:5
											localparam GPID_WIDTH = 1;
											// Trace: src/VX_gather_unit.sv:17:5
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam DATAW = 174;
											// Trace: src/VX_gather_unit.sv:18:5
											localparam DATA_WIS_OFF = 171;
											// Trace: src/VX_gather_unit.sv:19:5
											wire [0:0] result_in_valid;
											// Trace: src/VX_gather_unit.sv:20:5
											wire [173:0] result_in_data;
											// Trace: src/VX_gather_unit.sv:21:5
											wire [0:0] result_in_ready;
											// Trace: src/VX_gather_unit.sv:22:5
											localparam VX_gpu_pkg_ISSUE_ISW_BITS = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											wire [0:0] result_in_isw;
											// Trace: src/VX_gather_unit.sv:23:5
											genvar _gv_i_60;
											for (_gv_i_60 = 0; _gv_i_60 < BLOCK_SIZE; _gv_i_60 = _gv_i_60 + 1) begin : g_commit_in
												localparam i = _gv_i_60;
												// Trace: src/VX_gather_unit.sv:24:9
												assign result_in_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_result_if[i + _mbase_result_if].valid;
												// Trace: src/VX_gather_unit.sv:25:9
												assign result_in_data[i * 174+:174] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_result_if[i + _mbase_result_if].data;
												// Trace: src/VX_gather_unit.sv:26:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.lsu_unit.per_block_result_if[i + _mbase_result_if].ready = result_in_ready[i];
												if (1) begin : g_result_in_isw_full
													// Trace: src/VX_gather_unit.sv:34:13
													assign result_in_isw[i+:1] = sv2v_cast_1_signed(i);
												end
											end
											// Trace: src/VX_gather_unit.sv:37:5
											reg [0:0] result_out_valid;
											// Trace: src/VX_gather_unit.sv:38:5
											reg [173:0] result_out_data;
											// Trace: src/VX_gather_unit.sv:39:5
											wire [0:0] result_out_ready;
											// Trace: src/VX_gather_unit.sv:40:5
											always @(*) begin
												// Trace: src/VX_gather_unit.sv:41:9
												result_out_valid = 1'sb0;
												// Trace: src/VX_gather_unit.sv:42:9
												begin : sv2v_autoblock_12
													// Trace: src/VX_gather_unit.sv:42:14
													integer i;
													// Trace: src/VX_gather_unit.sv:42:14
													for (i = 0; i < 1; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:43:13
															result_out_data[i * 174+:174] = 1'sbx;
														end
												end
												begin : sv2v_autoblock_13
													// Trace: src/VX_gather_unit.sv:45:14
													integer i;
													// Trace: src/VX_gather_unit.sv:45:14
													for (i = 0; i < BLOCK_SIZE; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:46:13
															result_out_valid[result_in_isw[i+:1]] = result_in_valid[i];
															// Trace: src/VX_gather_unit.sv:47:13
															result_out_data[result_in_isw[i+:1] * 174+:174] = result_in_data[i * 174+:174];
														end
												end
											end
											// Trace: src/VX_gather_unit.sv:50:5
											genvar _gv_i_61;
											for (_gv_i_61 = 0; _gv_i_61 < BLOCK_SIZE; _gv_i_61 = _gv_i_61 + 1) begin : g_result_in_ready
												localparam i = _gv_i_61;
												// Trace: src/VX_gather_unit.sv:51:9
												assign result_in_ready[i] = result_out_ready[result_in_isw[i+:1]];
											end
											// Trace: src/VX_gather_unit.sv:53:5
											genvar _gv_i_62;
											localparam VX_gpu_pkg_SIMD_COUNT = 1;
											localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
											localparam VX_gpu_pkg_SIMD_IDX_W = 1;
											for (_gv_i_62 = 0; _gv_i_62 < 1; _gv_i_62 = _gv_i_62 + 1) begin : g_out_bufs
												localparam i = _gv_i_62;
												// Trace: src/VX_gather_unit.sv:54:9
												// expanded interface instance: result_tmp_if
												localparam _param_D4A7C_NUM_LANES = NUM_LANES;
												if (1) begin : result_tmp_if
													// removed import VX_gpu_pkg::*;
													// Trace: src/VX_result_if.sv:2:15
													localparam NUM_LANES = _param_D4A7C_NUM_LANES;
													// Trace: src/VX_result_if.sv:3:15
													localparam PID_WIDTH = 1;
													// Trace: src/VX_result_if.sv:5:5
													localparam VX_gpu_pkg_REG_TYPES = 1;
													localparam VX_gpu_pkg_RV_REGS = 32;
													localparam VX_gpu_pkg_NUM_REGS = 32;
													localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
													localparam VX_gpu_pkg_NW_BITS = 2;
													localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
													localparam VX_gpu_pkg_PC_BITS = 30;
													localparam VX_gpu_pkg_UUID_WIDTH = 1;
													// removed localparam type data_t
													// Trace: src/VX_result_if.sv:17:5
													wire valid;
													// Trace: src/VX_result_if.sv:18:5
													wire [173:0] data;
													// Trace: src/VX_result_if.sv:19:5
													wire ready;
													// Trace: src/VX_result_if.sv:20:5
													// Trace: src/VX_result_if.sv:25:5
												end
												// Trace: src/VX_gather_unit.sv:57:9
												VX_elastic_buffer #(
													.DATAW(DATAW),
													.SIZE(2),
													.OUT_REG(1)
												) out_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(result_out_valid[i]),
													.ready_in(result_out_ready[i]),
													.data_in(result_out_data[i * 174+:174]),
													.data_out(result_tmp_if.data),
													.valid_out(result_tmp_if.valid),
													.ready_out(result_tmp_if.ready)
												);
												// Trace: src/VX_gather_unit.sv:71:9
												wire [0:0] commit_sid_w;
												// Trace: src/VX_gather_unit.sv:72:9
												wire [3:0] commit_tmask_w;
												// Trace: src/VX_gather_unit.sv:73:9
												wire [127:0] commit_data_w;
												if (1) begin : g_no_lpid
													// Trace: src/VX_gather_unit.sv:91:13
													assign commit_sid_w = result_tmp_if.data[2];
													// Trace: src/VX_gather_unit.sv:92:13
													assign commit_tmask_w = result_tmp_if.data[170-:4];
													// Trace: src/VX_gather_unit.sv:93:13
													assign commit_data_w = result_tmp_if.data[130-:128];
												end
												// Trace: src/VX_gather_unit.sv:95:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_if].valid = result_tmp_if.valid;
												// Trace: src/VX_gather_unit.sv:96:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_if].data = {result_tmp_if.data[173], result_tmp_if.data[172-:2], commit_sid_w, commit_tmask_w, result_tmp_if.data[166-:30], result_tmp_if.data[136], result_tmp_if.data[135-:5], commit_data_w, result_tmp_if.data[1], result_tmp_if.data[0]};
												// Trace: src/VX_gather_unit.sv:108:9
												assign result_tmp_if.ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_if].ready;
											end
										end
										assign gather_unit.clk = clk;
										assign gather_unit.reset = reset;
									end
									assign lsu_unit.clk = clk;
									assign lsu_unit.reset = reset;
									// Trace: src/VX_execute.sv:35:5
									// expanded module instance: sfu_unit
									localparam _bbase_6660E_dispatch_if = 2;
									localparam _bbase_6660E_commit_if = 2;
									localparam _param_6660E_INSTANCE_ID = "";
									localparam _param_6660E_CORE_ID = CORE_ID;
									if (1) begin : sfu_unit
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_sfu_unit.sv:2:15
										localparam INSTANCE_ID = _param_6660E_INSTANCE_ID;
										// Trace: src/VX_sfu_unit.sv:3:15
										localparam CORE_ID = _param_6660E_CORE_ID;
										// Trace: src/VX_sfu_unit.sv:5:5
										wire clk;
										// Trace: src/VX_sfu_unit.sv:6:5
										wire reset;
										// Trace: src/VX_sfu_unit.sv:7:5
										// removed localparam type VX_gpu_pkg_base_dcrs_t
										wire [71:0] base_dcrs;
										// Trace: src/VX_sfu_unit.sv:8:5
										localparam _mbase_dispatch_if = 2;
										// Trace: src/VX_sfu_unit.sv:9:5
										// removed modport instance commit_csr_if
										// Trace: src/VX_sfu_unit.sv:10:5
										// removed modport instance sched_csr_if
										// Trace: src/VX_sfu_unit.sv:11:5
										localparam _mbase_commit_if = 2;
										// Trace: src/VX_sfu_unit.sv:12:5
										// removed modport instance warp_ctl_if
										// Trace: src/VX_sfu_unit.sv:14:5
										localparam BLOCK_SIZE = 1;
										// Trace: src/VX_sfu_unit.sv:15:5
										localparam NUM_LANES = 4;
										// Trace: src/VX_sfu_unit.sv:16:5
										localparam PE_COUNT = 2;
										// Trace: src/VX_sfu_unit.sv:17:5
										localparam PE_SEL_BITS = 1;
										// Trace: src/VX_sfu_unit.sv:18:5
										localparam PE_IDX_WCTL = 0;
										// Trace: src/VX_sfu_unit.sv:19:5
										localparam PE_IDX_CSRS = 1;
										// Trace: src/VX_sfu_unit.sv:20:5
										// expanded interface instance: per_block_execute_if
										localparam _param_E2592_NUM_LANES = NUM_LANES;
										genvar _arr_E2592;
										for (_arr_E2592 = 0; _arr_E2592 <= 0; _arr_E2592 = _arr_E2592 + 1) begin : per_block_execute_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_execute_if.sv:2:15
											localparam NUM_LANES = _param_E2592_NUM_LANES;
											// Trace: src/VX_execute_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_execute_if.sv:5:5
											localparam VX_gpu_pkg_INST_ALU_BITS = 4;
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
											// removed localparam type VX_gpu_pkg_alu_args_t
											localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
											// removed localparam type VX_gpu_pkg_csr_args_t
											localparam VX_gpu_pkg_INST_FMT_BITS = 2;
											localparam VX_gpu_pkg_INST_FRM_BITS = 3;
											// removed localparam type VX_gpu_pkg_fpu_args_t
											localparam VX_gpu_pkg_OFFSET_BITS = 12;
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											// removed localparam type data_t
											// Trace: src/VX_execute_if.sv:21:5
											wire valid;
											// Trace: src/VX_execute_if.sv:22:5
											wire [470:0] data;
											// Trace: src/VX_execute_if.sv:23:5
											wire ready;
											// Trace: src/VX_execute_if.sv:24:5
											// Trace: src/VX_execute_if.sv:29:5
										end
										// Trace: src/VX_sfu_unit.sv:23:5
										// expanded interface instance: per_block_result_if
										localparam _param_911F6_NUM_LANES = NUM_LANES;
										genvar _arr_911F6;
										for (_arr_911F6 = 0; _arr_911F6 <= 0; _arr_911F6 = _arr_911F6 + 1) begin : per_block_result_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_result_if.sv:2:15
											localparam NUM_LANES = _param_911F6_NUM_LANES;
											// Trace: src/VX_result_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_result_if.sv:5:5
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											// removed localparam type data_t
											// Trace: src/VX_result_if.sv:17:5
											wire valid;
											// Trace: src/VX_result_if.sv:18:5
											wire [173:0] data;
											// Trace: src/VX_result_if.sv:19:5
											wire ready;
											// Trace: src/VX_result_if.sv:20:5
											// Trace: src/VX_result_if.sv:25:5
										end
										// Trace: src/VX_sfu_unit.sv:26:5
										// expanded module instance: dispatch_unit
										localparam _bbase_2E16E_dispatch_if = 2;
										localparam _bbase_2E16E_execute_if = 0;
										localparam _param_2E16E_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_2E16E_NUM_LANES = NUM_LANES;
										localparam _param_2E16E_OUT_BUF = 3;
										if (1) begin : dispatch_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_dispatch_unit.sv:2:15
											localparam BLOCK_SIZE = _param_2E16E_BLOCK_SIZE;
											// Trace: src/VX_dispatch_unit.sv:3:15
											localparam NUM_LANES = _param_2E16E_NUM_LANES;
											// Trace: src/VX_dispatch_unit.sv:4:15
											localparam OUT_BUF = _param_2E16E_OUT_BUF;
											// Trace: src/VX_dispatch_unit.sv:5:15
											localparam MAX_FANOUT = 8;
											// Trace: src/VX_dispatch_unit.sv:7:5
											wire clk;
											// Trace: src/VX_dispatch_unit.sv:8:5
											wire reset;
											// Trace: src/VX_dispatch_unit.sv:9:5
											localparam _mbase_dispatch_if = 2;
											// Trace: src/VX_dispatch_unit.sv:10:5
											localparam _mbase_execute_if = 0;
											// Trace: src/VX_dispatch_unit.sv:12:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:13:5
											localparam NUM_PACKETS = 1;
											// Trace: src/VX_dispatch_unit.sv:14:5
											localparam LPID_BITS = 0;
											// Trace: src/VX_dispatch_unit.sv:15:5
											localparam LPID_WIDTH = 1;
											// Trace: src/VX_dispatch_unit.sv:16:5
											localparam GPID_BITS = 0;
											// Trace: src/VX_dispatch_unit.sv:17:5
											localparam GPID_WIDTH = 1;
											// Trace: src/VX_dispatch_unit.sv:18:5
											localparam BATCH_COUNT = 1;
											// Trace: src/VX_dispatch_unit.sv:19:5
											localparam BATCH_COUNT_W = 1;
											// Trace: src/VX_dispatch_unit.sv:20:5
											localparam ISSUE_W = 1;
											// Trace: src/VX_dispatch_unit.sv:21:5
											localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
											localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
											localparam VX_gpu_pkg_INST_OP_BITS = 4;
											localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
											localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
											localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NUM_SRC_OPDS = 3;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_SIMD_COUNT = 1;
											localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
											localparam VX_gpu_pkg_SIMD_IDX_W = 1;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam IN_DATAW = 471;
											// Trace: src/VX_dispatch_unit.sv:22:5
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam OUT_DATAW = 471;
											// Trace: src/VX_dispatch_unit.sv:23:5
											localparam FANOUT_ENABLE = 1'd0;
											// Trace: src/VX_dispatch_unit.sv:24:5
											localparam DATA_TMASK_OFF = 463;
											// Trace: src/VX_dispatch_unit.sv:25:5
											localparam DATA_REGS_OFF = 2;
											// Trace: src/VX_dispatch_unit.sv:26:5
											// removed localparam type packet_t
											// Trace: src/VX_dispatch_unit.sv:30:5
											wire [0:0] dispatch_valid;
											// Trace: src/VX_dispatch_unit.sv:31:5
											wire [470:0] dispatch_data;
											// Trace: src/VX_dispatch_unit.sv:32:5
											wire [0:0] dispatch_ready;
											// Trace: src/VX_dispatch_unit.sv:33:5
											genvar _gv_i_35;
											for (_gv_i_35 = 0; _gv_i_35 < 1; _gv_i_35 = _gv_i_35 + 1) begin : g_dispatch_data
												localparam i = _gv_i_35;
												// Trace: src/VX_dispatch_unit.sv:34:9
												assign dispatch_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].valid;
												// Trace: src/VX_dispatch_unit.sv:35:9
												assign dispatch_data[i * 471+:471] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].data;
												// Trace: src/VX_dispatch_unit.sv:36:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.dispatch_if[i + _mbase_dispatch_if].ready = dispatch_ready[i];
											end
											// Trace: src/VX_dispatch_unit.sv:38:5
											wire [0:0] block_ready;
											// Trace: src/VX_dispatch_unit.sv:39:5
											wire [3:0] block_tmask;
											// Trace: src/VX_dispatch_unit.sv:40:5
											wire [383:0] block_rsdata;
											// Trace: src/VX_dispatch_unit.sv:41:5
											wire [0:0] block_pid;
											// Trace: src/VX_dispatch_unit.sv:42:5
											wire [0:0] block_sop;
											// Trace: src/VX_dispatch_unit.sv:43:5
											wire [0:0] block_eop;
											// Trace: src/VX_dispatch_unit.sv:44:5
											wire [0:0] block_done;
											// Trace: src/VX_dispatch_unit.sv:45:5
											wire batch_done = &block_done;
											// Trace: src/VX_dispatch_unit.sv:46:5
											wire [0:0] batch_idx;
											// Trace: src/VX_dispatch_unit.sv:47:5
											if (1) begin : g_batch_idx_0
												// Trace: src/VX_dispatch_unit.sv:73:9
												assign batch_idx = 0;
											end
											// Trace: src/VX_dispatch_unit.sv:75:5
											wire [0:0] issue_indices;
											// Trace: src/VX_dispatch_unit.sv:76:5
											genvar _gv_block_idx_2;
											for (_gv_block_idx_2 = 0; _gv_block_idx_2 < BLOCK_SIZE; _gv_block_idx_2 = _gv_block_idx_2 + 1) begin : g_issue_indices
												localparam block_idx = _gv_block_idx_2;
												// Trace: src/VX_dispatch_unit.sv:77:9
												assign issue_indices[block_idx+:1] = sv2v_cast_1(batch_idx * BLOCK_SIZE) + sv2v_cast_1_signed(block_idx);
											end
											// Trace: src/VX_dispatch_unit.sv:79:5
											genvar _gv_block_idx_3;
											localparam VX_gpu_pkg_ISSUE_ISW_BITS = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											function automatic [1:0] VX_gpu_pkg_wis_to_wid;
												// Trace: src/VX_gpu_pkg.sv:264:9
												input reg [1:0] wis;
												// Trace: src/VX_gpu_pkg.sv:265:9
												input reg [0:0] isw;
												// Trace: src/VX_gpu_pkg.sv:267:9
												begin
													// Trace: src/VX_gpu_pkg.sv:270:13
													VX_gpu_pkg_wis_to_wid = wis;
												end
											endfunction
											for (_gv_block_idx_3 = 0; _gv_block_idx_3 < BLOCK_SIZE; _gv_block_idx_3 = _gv_block_idx_3 + 1) begin : g_blocks
												localparam block_idx = _gv_block_idx_3;
												// Trace: src/VX_dispatch_unit.sv:80:9
												wire [0:0] issue_idx = issue_indices[block_idx+:1];
												// Trace: src/VX_dispatch_unit.sv:81:9
												wire [1:0] dispatch_wis = dispatch_data[(issue_idx * 471) + 468+:VX_gpu_pkg_ISSUE_WIS_W];
												// Trace: src/VX_dispatch_unit.sv:82:9
												wire [0:0] dispatch_sid = dispatch_data[(issue_idx * 471) + 467+:VX_gpu_pkg_SIMD_IDX_W];
												// Trace: src/VX_dispatch_unit.sv:83:9
												wire dispatch_sop = dispatch_data[(issue_idx * 471) + 1];
												// Trace: src/VX_dispatch_unit.sv:84:9
												wire dispatch_eop = dispatch_data[issue_idx * 471];
												// Trace: src/VX_dispatch_unit.sv:85:9
												wire [3:0] dispatch_tmask;
												// Trace: src/VX_dispatch_unit.sv:86:9
												wire [383:0] dispatch_rsdata;
												// Trace: src/VX_dispatch_unit.sv:87:9
												assign dispatch_tmask = dispatch_data[(issue_idx * 471) + DATA_TMASK_OFF+:4];
												// Trace: src/VX_dispatch_unit.sv:88:9
												assign dispatch_rsdata[0+:128] = dispatch_data[(issue_idx * 471) + 258+:128];
												// Trace: src/VX_dispatch_unit.sv:89:9
												assign dispatch_rsdata[128+:128] = dispatch_data[(issue_idx * 471) + 130+:128];
												// Trace: src/VX_dispatch_unit.sv:90:9
												assign dispatch_rsdata[256+:128] = dispatch_data[(issue_idx * 471) + 2+:128];
												// Trace: src/VX_dispatch_unit.sv:91:9
												wire valid_p;
												wire ready_p;
												if (1) begin : g_full_simd
													// Trace: src/VX_dispatch_unit.sv:132:13
													assign valid_p = dispatch_valid[issue_idx];
													// Trace: src/VX_dispatch_unit.sv:133:13
													assign block_tmask[block_idx * 4+:4] = dispatch_tmask;
													// Trace: src/VX_dispatch_unit.sv:134:13
													assign block_rsdata[32 * (4 * (block_idx * 3))+:384] = dispatch_rsdata;
													// Trace: src/VX_dispatch_unit.sv:135:13
													assign block_pid[block_idx+:1] = 0;
													// Trace: src/VX_dispatch_unit.sv:136:13
													assign block_sop[block_idx] = 1;
													// Trace: src/VX_dispatch_unit.sv:137:13
													assign block_eop[block_idx] = 1;
													// Trace: src/VX_dispatch_unit.sv:138:13
													assign block_ready[block_idx] = ready_p;
													// Trace: src/VX_dispatch_unit.sv:139:13
													assign block_done[block_idx] = ready_p || ~valid_p;
												end
												// Trace: src/VX_dispatch_unit.sv:141:9
												wire [0:0] isw;
												if (1) begin : g_isw
													// Trace: src/VX_dispatch_unit.sv:149:13
													assign isw = block_idx;
												end
												// Trace: src/VX_dispatch_unit.sv:151:9
												wire [1:0] block_wid = VX_gpu_pkg_wis_to_wid(dispatch_wis, isw);
												// Trace: src/VX_dispatch_unit.sv:152:9
												wire [0:0] warp_pid = block_pid[block_idx+:1] + sv2v_cast_1(dispatch_sid * NUM_PACKETS);
												// Trace: src/VX_dispatch_unit.sv:153:9
												wire warp_sop = block_sop[block_idx] && dispatch_sop;
												// Trace: src/VX_dispatch_unit.sv:154:9
												wire warp_eop = block_eop[block_idx] && dispatch_eop;
												// Trace: src/VX_dispatch_unit.sv:155:9
												VX_elastic_buffer #(
													.DATAW(OUT_DATAW),
													.SIZE(2),
													.OUT_REG(1)
												) buf_out(
													.clk(clk),
													.reset(reset),
													.valid_in(valid_p),
													.ready_in(ready_p),
													.data_in({dispatch_data[(issue_idx * 471) + 470-:VX_gpu_pkg_UUID_WIDTH], block_wid, block_tmask[block_idx * 4+:4], dispatch_data[(issue_idx * 471) + 462-:77], block_rsdata[32 * ((block_idx * 3) * 4)+:128], block_rsdata[32 * (((block_idx * 3) + 1) * 4)+:128], block_rsdata[32 * (((block_idx * 3) + 2) * 4)+:128], warp_pid, warp_sop, warp_eop}),
													.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_execute_if[block_idx + _mbase_execute_if].data),
													.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_execute_if[block_idx + _mbase_execute_if].valid),
													.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_execute_if[block_idx + _mbase_execute_if].ready)
												);
											end
											// Trace: src/VX_dispatch_unit.sv:180:5
											reg [0:0] ready_in;
											// Trace: src/VX_dispatch_unit.sv:181:5
											always @(*) begin
												// Trace: src/VX_dispatch_unit.sv:182:9
												ready_in = 0;
												// Trace: src/VX_dispatch_unit.sv:183:9
												begin : sv2v_autoblock_14
													// Trace: src/VX_dispatch_unit.sv:183:14
													integer block_idx;
													// Trace: src/VX_dispatch_unit.sv:183:14
													for (block_idx = 0; block_idx < BLOCK_SIZE; block_idx = block_idx + 1)
														begin
															// Trace: src/VX_dispatch_unit.sv:184:13
															ready_in[issue_indices[block_idx+:1]] = block_ready[block_idx] && block_eop[block_idx];
														end
												end
											end
											// Trace: src/VX_dispatch_unit.sv:187:5
											assign dispatch_ready = ready_in;
										end
										assign dispatch_unit.clk = clk;
										assign dispatch_unit.reset = reset;
										// Trace: src/VX_sfu_unit.sv:36:5
										// expanded interface instance: pe_execute_if
										localparam _param_C9035_NUM_LANES = NUM_LANES;
										genvar _arr_C9035;
										for (_arr_C9035 = 0; _arr_C9035 <= 1; _arr_C9035 = _arr_C9035 + 1) begin : pe_execute_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_execute_if.sv:2:15
											localparam NUM_LANES = _param_C9035_NUM_LANES;
											// Trace: src/VX_execute_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_execute_if.sv:5:5
											localparam VX_gpu_pkg_INST_ALU_BITS = 4;
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
											// removed localparam type VX_gpu_pkg_alu_args_t
											localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
											// removed localparam type VX_gpu_pkg_csr_args_t
											localparam VX_gpu_pkg_INST_FMT_BITS = 2;
											localparam VX_gpu_pkg_INST_FRM_BITS = 3;
											// removed localparam type VX_gpu_pkg_fpu_args_t
											localparam VX_gpu_pkg_OFFSET_BITS = 12;
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											// removed localparam type data_t
											// Trace: src/VX_execute_if.sv:21:5
											wire valid;
											// Trace: src/VX_execute_if.sv:22:5
											wire [470:0] data;
											// Trace: src/VX_execute_if.sv:23:5
											wire ready;
											// Trace: src/VX_execute_if.sv:24:5
											// Trace: src/VX_execute_if.sv:29:5
										end
										// Trace: src/VX_sfu_unit.sv:39:5
										// expanded interface instance: pe_result_if
										localparam _param_FE18D_NUM_LANES = NUM_LANES;
										genvar _arr_FE18D;
										for (_arr_FE18D = 0; _arr_FE18D <= 1; _arr_FE18D = _arr_FE18D + 1) begin : pe_result_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_result_if.sv:2:15
											localparam NUM_LANES = _param_FE18D_NUM_LANES;
											// Trace: src/VX_result_if.sv:3:15
											localparam PID_WIDTH = 1;
											// Trace: src/VX_result_if.sv:5:5
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											// removed localparam type data_t
											// Trace: src/VX_result_if.sv:17:5
											wire valid;
											// Trace: src/VX_result_if.sv:18:5
											wire [173:0] data;
											// Trace: src/VX_result_if.sv:19:5
											wire ready;
											// Trace: src/VX_result_if.sv:20:5
											// Trace: src/VX_result_if.sv:25:5
										end
										// Trace: src/VX_sfu_unit.sv:42:5
										reg [0:0] pe_select;
										// Trace: src/VX_sfu_unit.sv:43:5
										localparam VX_gpu_pkg_INST_SFU_BITS = 4;
										function automatic VX_gpu_pkg_inst_sfu_is_csr;
											// Trace: src/VX_gpu_pkg.sv:255:46
											input reg [3:0] op;
											// Trace: src/VX_gpu_pkg.sv:256:9
											VX_gpu_pkg_inst_sfu_is_csr = (op >= 6) && (op <= 8);
										endfunction
										always @(*) begin
											// Trace: src/VX_sfu_unit.sv:44:9
											pe_select = PE_IDX_WCTL;
											// Trace: src/VX_sfu_unit.sv:45:9
											if (VX_gpu_pkg_inst_sfu_is_csr(per_block_execute_if[0].data[433-:4]))
												// Trace: src/VX_sfu_unit.sv:46:13
												pe_select = PE_IDX_CSRS;
										end
										// Trace: src/VX_sfu_unit.sv:49:5
										// expanded module instance: pe_switch
										localparam _bbase_3D12E_execute_in_if = 0;
										localparam _bbase_3D12E_result_out_if = 0;
										localparam _bbase_3D12E_execute_out_if = 0;
										localparam _bbase_3D12E_result_in_if = 0;
										localparam _param_3D12E_PE_COUNT = PE_COUNT;
										localparam _param_3D12E_NUM_LANES = NUM_LANES;
										localparam _param_3D12E_ARBITER = "R";
										localparam _param_3D12E_REQ_OUT_BUF = 0;
										localparam _param_3D12E_RSP_OUT_BUF = 3;
										if (1) begin : pe_switch
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_pe_switch.sv:2:15
											localparam PE_COUNT = _param_3D12E_PE_COUNT;
											// Trace: src/VX_pe_switch.sv:3:15
											localparam NUM_LANES = _param_3D12E_NUM_LANES;
											// Trace: src/VX_pe_switch.sv:4:15
											localparam REQ_OUT_BUF = _param_3D12E_REQ_OUT_BUF;
											// Trace: src/VX_pe_switch.sv:5:15
											localparam RSP_OUT_BUF = _param_3D12E_RSP_OUT_BUF;
											// Trace: src/VX_pe_switch.sv:6:15
											localparam ARBITER = _param_3D12E_ARBITER;
											// Trace: src/VX_pe_switch.sv:7:15
											localparam PE_SEL_BITS = 1;
											// Trace: src/VX_pe_switch.sv:9:5
											wire clk;
											// Trace: src/VX_pe_switch.sv:10:5
											wire reset;
											// Trace: src/VX_pe_switch.sv:11:5
											wire [0:0] pe_sel;
											// Trace: src/VX_pe_switch.sv:12:5
											localparam _mbase_execute_in_if = _bbase_3D12E_execute_in_if;
											// Trace: src/VX_pe_switch.sv:13:5
											localparam _mbase_result_out_if = _bbase_3D12E_result_out_if;
											// Trace: src/VX_pe_switch.sv:14:5
											localparam _mbase_execute_out_if = 0;
											// Trace: src/VX_pe_switch.sv:15:5
											localparam _mbase_result_in_if = 0;
											// Trace: src/VX_pe_switch.sv:17:5
											localparam PID_BITS = 0;
											// Trace: src/VX_pe_switch.sv:18:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_pe_switch.sv:19:5
											localparam VX_gpu_pkg_INST_ALU_BITS = 4;
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam VX_gpu_pkg_ALU_TYPE_BITS = 2;
											// removed localparam type VX_gpu_pkg_alu_args_t
											localparam VX_gpu_pkg_INST_ARGS_BITS = 37;
											// removed localparam type VX_gpu_pkg_csr_args_t
											localparam VX_gpu_pkg_INST_FMT_BITS = 2;
											localparam VX_gpu_pkg_INST_FRM_BITS = 3;
											// removed localparam type VX_gpu_pkg_fpu_args_t
											localparam VX_gpu_pkg_OFFSET_BITS = 12;
											// removed localparam type VX_gpu_pkg_lsu_args_t
											// removed localparam type VX_gpu_pkg_wctl_args_t
											// removed localparam type VX_gpu_pkg_op_args_t
											localparam REQ_DATAW = 471;
											// Trace: src/VX_pe_switch.sv:20:5
											localparam RSP_DATAW = 174;
											// Trace: src/VX_pe_switch.sv:21:5
											wire [1:0] pe_req_valid;
											// Trace: src/VX_pe_switch.sv:22:5
											wire [941:0] pe_req_data;
											// Trace: src/VX_pe_switch.sv:23:5
											wire [1:0] pe_req_ready;
											// Trace: src/VX_pe_switch.sv:24:5
											VX_stream_switch #(
												.DATAW(REQ_DATAW),
												.NUM_INPUTS(1),
												.NUM_OUTPUTS(PE_COUNT),
												.OUT_BUF(REQ_OUT_BUF)
											) req_switch(
												.clk(clk),
												.reset(reset),
												.sel_in(pe_sel),
												.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_execute_if[_mbase_execute_in_if].valid),
												.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_execute_if[_mbase_execute_in_if].ready),
												.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_execute_if[_mbase_execute_in_if].data),
												.data_out(pe_req_data),
												.valid_out(pe_req_valid),
												.ready_out(pe_req_ready)
											);
											// Trace: src/VX_pe_switch.sv:40:5
											genvar _gv_i_150;
											for (_gv_i_150 = 0; _gv_i_150 < PE_COUNT; _gv_i_150 = _gv_i_150 + 1) begin : g_execute_out_if
												localparam i = _gv_i_150;
												// Trace: src/VX_pe_switch.sv:41:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[i + _mbase_execute_out_if].valid = pe_req_valid[i];
												// Trace: src/VX_pe_switch.sv:42:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[i + _mbase_execute_out_if].data = pe_req_data[i * 471+:471];
												// Trace: src/VX_pe_switch.sv:43:9
												assign pe_req_ready[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[i + _mbase_execute_out_if].ready;
											end
											// Trace: src/VX_pe_switch.sv:45:5
											wire [1:0] pe_rsp_valid;
											// Trace: src/VX_pe_switch.sv:46:5
											wire [347:0] pe_rsp_data;
											// Trace: src/VX_pe_switch.sv:47:5
											wire [1:0] pe_rsp_ready;
											// Trace: src/VX_pe_switch.sv:48:5
											genvar _gv_i_151;
											for (_gv_i_151 = 0; _gv_i_151 < PE_COUNT; _gv_i_151 = _gv_i_151 + 1) begin : g_result_in_if
												localparam i = _gv_i_151;
												// Trace: src/VX_pe_switch.sv:49:9
												assign pe_rsp_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[i + _mbase_result_in_if].valid;
												// Trace: src/VX_pe_switch.sv:50:9
												assign pe_rsp_data[i * 174+:174] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[i + _mbase_result_in_if].data;
												// Trace: src/VX_pe_switch.sv:51:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[i + _mbase_result_in_if].ready = pe_rsp_ready[i];
											end
											// Trace: src/VX_pe_switch.sv:53:5
											VX_stream_arb #(
												.NUM_INPUTS(PE_COUNT),
												.DATAW(RSP_DATAW),
												.ARBITER(ARBITER),
												.OUT_BUF(RSP_OUT_BUF)
											) rsp_arb(
												.clk(clk),
												.reset(reset),
												.valid_in(pe_rsp_valid),
												.ready_in(pe_rsp_ready),
												.data_in(pe_rsp_data),
												.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_result_if[_mbase_result_out_if].data),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_result_if[_mbase_result_out_if].valid),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_result_if[_mbase_result_out_if].ready),
												.sel_out()
											);
										end
										assign pe_switch.clk = clk;
										assign pe_switch.reset = reset;
										assign pe_switch.pe_sel = pe_select;
										// Trace: src/VX_sfu_unit.sv:64:5
										// expanded module instance: wctl_unit
										localparam _bbase_F22EA_execute_if = PE_IDX_WCTL;
										localparam _bbase_F22EA_result_if = PE_IDX_WCTL;
										localparam _param_F22EA_INSTANCE_ID = "";
										localparam _param_F22EA_NUM_LANES = NUM_LANES;
										if (1) begin : wctl_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_wctl_unit.sv:2:15
											localparam INSTANCE_ID = _param_F22EA_INSTANCE_ID;
											// Trace: src/VX_wctl_unit.sv:3:15
											localparam NUM_LANES = _param_F22EA_NUM_LANES;
											// Trace: src/VX_wctl_unit.sv:5:5
											wire clk;
											// Trace: src/VX_wctl_unit.sv:6:5
											wire reset;
											// Trace: src/VX_wctl_unit.sv:7:5
											localparam _mbase_execute_if = _bbase_F22EA_execute_if;
											// Trace: src/VX_wctl_unit.sv:8:5
											// removed modport instance warp_ctl_if
											// Trace: src/VX_wctl_unit.sv:9:5
											localparam _mbase_result_if = _bbase_F22EA_result_if;
											// Trace: src/VX_wctl_unit.sv:11:5
											localparam LANE_BITS = 2;
											// Trace: src/VX_wctl_unit.sv:12:5
											localparam PID_BITS = 0;
											// Trace: src/VX_wctl_unit.sv:13:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_wctl_unit.sv:14:5
											localparam VX_gpu_pkg_NB_BITS = 1;
											localparam VX_gpu_pkg_NB_WIDTH = VX_gpu_pkg_NB_BITS;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											// removed localparam type VX_gpu_pkg_barrier_t
											localparam VX_gpu_pkg_DV_STACK_SIZE = 3;
											localparam VX_gpu_pkg_DV_STACK_SIZEW = 2;
											// removed localparam type VX_gpu_pkg_join_t
											localparam VX_gpu_pkg_PC_BITS = 30;
											// removed localparam type VX_gpu_pkg_split_t
											// removed localparam type VX_gpu_pkg_tmc_t
											// removed localparam type VX_gpu_pkg_wspawn_t
											localparam WCTL_WIDTH = 89;
											// Trace: src/VX_wctl_unit.sv:15:5
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam DATAW = 48;
											// Trace: src/VX_wctl_unit.sv:16:5
											wire [4:0] tmc;
											// Trace: src/VX_wctl_unit.sv:17:5
											wire [34:0] wspawn;
											// Trace: src/VX_wctl_unit.sv:18:5
											wire [39:0] split;
											// Trace: src/VX_wctl_unit.sv:19:5
											wire [2:0] sjoin;
											// Trace: src/VX_wctl_unit.sv:20:5
											wire [5:0] barrier;
											// Trace: src/VX_wctl_unit.sv:21:5
											localparam VX_gpu_pkg_INST_SFU_WSPAWN = 4'h1;
											wire is_wspawn = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[433-:4] == VX_gpu_pkg_INST_SFU_WSPAWN;
											// Trace: src/VX_wctl_unit.sv:22:5
											localparam VX_gpu_pkg_INST_SFU_TMC = 4'h0;
											wire is_tmc = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[433-:4] == VX_gpu_pkg_INST_SFU_TMC;
											// Trace: src/VX_wctl_unit.sv:23:5
											localparam VX_gpu_pkg_INST_SFU_PRED = 4'h5;
											wire is_pred = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[433-:4] == VX_gpu_pkg_INST_SFU_PRED;
											// Trace: src/VX_wctl_unit.sv:24:5
											localparam VX_gpu_pkg_INST_SFU_SPLIT = 4'h2;
											wire is_split = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[433-:4] == VX_gpu_pkg_INST_SFU_SPLIT;
											// Trace: src/VX_wctl_unit.sv:25:5
											localparam VX_gpu_pkg_INST_SFU_JOIN = 4'h3;
											wire is_join = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[433-:4] == VX_gpu_pkg_INST_SFU_JOIN;
											// Trace: src/VX_wctl_unit.sv:26:5
											localparam VX_gpu_pkg_INST_SFU_BAR = 4'h4;
											wire is_bar = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[433-:4] == VX_gpu_pkg_INST_SFU_BAR;
											// Trace: src/VX_wctl_unit.sv:27:5
											wire [1:0] last_tid;
											// Trace: src/VX_wctl_unit.sv:28:5
											if (1) begin : g_last_tid
												// Trace: src/VX_wctl_unit.sv:29:9
												VX_priority_encoder #(
													.N(NUM_LANES),
													.REVERSE(1)
												) last_tid_select(
													.data_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[467-:4]),
													.index_out(last_tid),
													.onehot_out(),
													.valid_out()
												);
											end
											// Trace: src/VX_wctl_unit.sv:41:5
											wire [31:0] rs1_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[259 + (last_tid * 32)+:32];
											// Trace: src/VX_wctl_unit.sv:42:5
											wire [31:0] rs2_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[131 + (last_tid * 32)+:32];
											// Trace: src/VX_wctl_unit.sv:43:5
											wire not_pred = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[393];
											// Trace: src/VX_wctl_unit.sv:44:5
											wire [3:0] taken;
											// Trace: src/VX_wctl_unit.sv:45:5
											genvar _gv_i_138;
											for (_gv_i_138 = 0; _gv_i_138 < NUM_LANES; _gv_i_138 = _gv_i_138 + 1) begin : g_taken
												localparam i = _gv_i_138;
												// Trace: src/VX_wctl_unit.sv:46:9
												assign taken[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[259 + (i * 32)] ^ not_pred;
											end
											// Trace: src/VX_wctl_unit.sv:48:5
											wire [3:0] then_tmask;
											// Trace: src/VX_wctl_unit.sv:49:5
											wire [3:0] else_tmask;
											// Trace: src/VX_wctl_unit.sv:50:5
											if (1) begin : g_no_pid
												// Trace: src/VX_wctl_unit.sv:64:9
												assign then_tmask = taken & Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[467-:4];
												// Trace: src/VX_wctl_unit.sv:65:9
												assign else_tmask = ~taken & Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[467-:4];
											end
											// Trace: src/VX_wctl_unit.sv:67:5
											wire has_then = then_tmask != 0;
											// Trace: src/VX_wctl_unit.sv:68:5
											wire has_else = else_tmask != 0;
											// Trace: src/VX_wctl_unit.sv:69:5
											wire [3:0] pred_mask = (has_then ? then_tmask : rs2_data[3:0]);
											// Trace: src/VX_wctl_unit.sv:70:5
											assign tmc[4] = is_tmc || is_pred;
											// Trace: src/VX_wctl_unit.sv:71:5
											assign tmc[3-:4] = (is_pred ? pred_mask : rs1_data[3:0]);
											// Trace: src/VX_wctl_unit.sv:72:5
											wire [2:0] then_tmask_cnt;
											wire [2:0] else_tmask_cnt;
											// Trace: src/VX_wctl_unit.sv:73:5
											VX_popcount #(
												.N(4),
												.MODEL(1)
											) __pop_count_ex114(
												.data_in(then_tmask),
												.data_out(then_tmask_cnt)
											);
											// Trace: src/VX_wctl_unit.sv:80:5
											VX_popcount #(
												.N(4),
												.MODEL(1)
											) __pop_count_ex115(
												.data_in(else_tmask),
												.data_out(else_tmask_cnt)
											);
											// Trace: src/VX_wctl_unit.sv:87:5
											wire then_first = then_tmask_cnt >= else_tmask_cnt;
											// Trace: src/VX_wctl_unit.sv:88:5
											wire [3:0] taken_tmask = (then_first ? then_tmask : else_tmask);
											// Trace: src/VX_wctl_unit.sv:89:5
											wire [3:0] ntaken_tmask = (then_first ? else_tmask : then_tmask);
											// Trace: src/VX_wctl_unit.sv:90:5
											assign split[39] = is_split;
											// Trace: src/VX_wctl_unit.sv:91:5
											assign split[38] = has_then && has_else;
											// Trace: src/VX_wctl_unit.sv:92:5
											assign split[37-:4] = taken_tmask;
											// Trace: src/VX_wctl_unit.sv:93:5
											assign split[33-:4] = ntaken_tmask;
											// Trace: src/VX_wctl_unit.sv:94:5
											function automatic [29:0] VX_gpu_pkg_from_fullPC;
												// Trace: src/VX_gpu_pkg.sv:30:56
												input reg [31:0] pc;
												// Trace: src/VX_gpu_pkg.sv:31:9
												VX_gpu_pkg_from_fullPC = sv2v_cast_30(pc >> 2);
											endfunction
											assign split[29-:30] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[463-:30] + VX_gpu_pkg_from_fullPC(32'sd4);
											// Trace: src/VX_wctl_unit.sv:95:5
											assign sjoin[2] = is_join;
											// Trace: src/VX_wctl_unit.sv:96:5
											assign sjoin[1-:2] = rs1_data[1:0];
											// Trace: src/VX_wctl_unit.sv:97:5
											assign barrier[5] = is_bar;
											// Trace: src/VX_wctl_unit.sv:98:5
											assign barrier[4-:1] = rs1_data[0:0];
											// Trace: src/VX_wctl_unit.sv:99:5
											assign barrier[3] = 1'b0;
											// Trace: src/VX_wctl_unit.sv:100:5
											function automatic signed [1:0] sv2v_cast_8835B_signed;
												input reg signed [1:0] inp;
												sv2v_cast_8835B_signed = inp;
											endfunction
											assign barrier[2-:2] = rs2_data[1:0] - sv2v_cast_8835B_signed(1);
											// Trace: src/VX_wctl_unit.sv:101:5
											assign barrier[0] = rs2_data[1:0] == sv2v_cast_8835B_signed(1);
											// Trace: src/VX_wctl_unit.sv:102:5
											wire [3:0] wspawn_wmask;
											// Trace: src/VX_wctl_unit.sv:103:5
											genvar _gv_i_139;
											for (_gv_i_139 = 0; _gv_i_139 < 4; _gv_i_139 = _gv_i_139 + 1) begin : g_wspawn_wmask
												localparam i = _gv_i_139;
												// Trace: src/VX_wctl_unit.sv:104:9
												assign wspawn_wmask[i] = (i < rs1_data[VX_gpu_pkg_NW_BITS:0]) && (i != Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[469-:2]);
											end
											// Trace: src/VX_wctl_unit.sv:106:5
											assign wspawn[34] = is_wspawn;
											// Trace: src/VX_wctl_unit.sv:107:5
											assign wspawn[33-:4] = wspawn_wmask;
											// Trace: src/VX_wctl_unit.sv:108:5
											assign wspawn[29-:30] = VX_gpu_pkg_from_fullPC(rs2_data);
											// Trace: src/VX_wctl_unit.sv:109:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.dvstack_wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[469-:2];
											// Trace: src/VX_wctl_unit.sv:110:5
											wire [1:0] dvstack_ptr;
											// Trace: src/VX_wctl_unit.sv:111:5
											VX_elastic_buffer #(
												.DATAW(DATAW),
												.SIZE(2)
											) rsp_buf(
												.clk(clk),
												.reset(reset),
												.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].valid),
												.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].ready),
												.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[470], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[469-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[467-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[463-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[391-:5], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[392], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[0], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.dvstack_ptr}),
												.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[173], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[172-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[170-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[166-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[135-:5], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[136], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[0], dvstack_ptr}),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].valid),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].ready)
											);
											// Trace: src/VX_wctl_unit.sv:124:5
											wire execute_fire = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].valid && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].ready;
											// Trace: src/VX_wctl_unit.sv:125:5
											wire wctl_valid = execute_fire && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[0];
											// Trace: src/VX_wctl_unit.sv:126:5
											VX_pipe_register #(
												.DATAW(92),
												.RESETW(1)
											) wctl_reg(
												.clk(clk),
												.reset(reset),
												.enable(1'b1),
												.data_in({wctl_valid, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[469-:2], tmc, wspawn, split, sjoin, barrier}),
												.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.valid, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wid, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.tmc, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.wspawn, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.split, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.sjoin, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.warp_ctl_if.barrier})
											);
											// Trace: src/VX_wctl_unit.sv:136:5
											genvar _gv_i_140;
											for (_gv_i_140 = 0; _gv_i_140 < NUM_LANES; _gv_i_140 = _gv_i_140 + 1) begin : g_result_if
												localparam i = _gv_i_140;
												// Trace: src/VX_wctl_unit.sv:137:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[3 + (i * 32)+:32] = sv2v_cast_32(dvstack_ptr);
											end
										end
										assign wctl_unit.clk = clk;
										assign wctl_unit.reset = reset;
										// Trace: src/VX_sfu_unit.sv:74:5
										// expanded module instance: csr_unit
										localparam _bbase_BED2E_execute_if = PE_IDX_CSRS;
										localparam _bbase_BED2E_result_if = PE_IDX_CSRS;
										localparam _param_BED2E_INSTANCE_ID = "";
										localparam _param_BED2E_CORE_ID = CORE_ID;
										localparam _param_BED2E_NUM_LANES = NUM_LANES;
										if (1) begin : csr_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_csr_unit.sv:2:15
											localparam INSTANCE_ID = _param_BED2E_INSTANCE_ID;
											// Trace: src/VX_csr_unit.sv:3:15
											localparam CORE_ID = _param_BED2E_CORE_ID;
											// Trace: src/VX_csr_unit.sv:4:15
											localparam NUM_LANES = _param_BED2E_NUM_LANES;
											// Trace: src/VX_csr_unit.sv:6:5
											wire clk;
											// Trace: src/VX_csr_unit.sv:7:5
											wire reset;
											// Trace: src/VX_csr_unit.sv:8:5
											// removed localparam type VX_gpu_pkg_base_dcrs_t
											wire [71:0] base_dcrs;
											// Trace: src/VX_csr_unit.sv:9:5
											// removed modport instance commit_csr_if
											// Trace: src/VX_csr_unit.sv:10:5
											// removed modport instance sched_csr_if
											// Trace: src/VX_csr_unit.sv:11:5
											localparam _mbase_execute_if = _bbase_BED2E_execute_if;
											// Trace: src/VX_csr_unit.sv:12:5
											localparam _mbase_result_if = _bbase_BED2E_result_if;
											// Trace: src/VX_csr_unit.sv:14:5
											localparam PID_BITS = 0;
											// Trace: src/VX_csr_unit.sv:15:5
											localparam PID_WIDTH = 1;
											// Trace: src/VX_csr_unit.sv:16:5
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam DATAW = 174;
											// Trace: src/VX_csr_unit.sv:17:5
											reg [127:0] csr_read_data;
											// Trace: src/VX_csr_unit.sv:18:5
											reg [31:0] csr_write_data;
											// Trace: src/VX_csr_unit.sv:19:5
											wire [31:0] csr_read_data_ro;
											wire [31:0] csr_read_data_rw;
											// Trace: src/VX_csr_unit.sv:20:5
											wire [31:0] csr_req_data;
											// Trace: src/VX_csr_unit.sv:21:5
											reg csr_rd_enable;
											// Trace: src/VX_csr_unit.sv:22:5
											wire csr_wr_enable;
											// Trace: src/VX_csr_unit.sv:23:5
											wire csr_req_ready;
											// Trace: src/VX_csr_unit.sv:24:5
											wire [11:0] csr_addr = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[409-:12];
											// Trace: src/VX_csr_unit.sv:25:5
											localparam VX_gpu_pkg_RV_REGS_BITS = 5;
											wire [4:0] csr_imm = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[397-:5];
											// Trace: src/VX_csr_unit.sv:26:5
											wire is_fpu_csr = csr_addr <= 12'h003;
											// Trace: src/VX_csr_unit.sv:27:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.alm_empty_wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[469-:2];
											// Trace: src/VX_csr_unit.sv:28:5
											wire no_pending_instr = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.alm_empty || ~is_fpu_csr;
											// Trace: src/VX_csr_unit.sv:29:5
											wire csr_req_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].valid && no_pending_instr;
											// Trace: src/VX_csr_unit.sv:30:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].ready = csr_req_ready && no_pending_instr;
											// Trace: src/VX_csr_unit.sv:31:5
											wire [127:0] rs1_data;
											// Trace: src/VX_csr_unit.sv:32:5
											genvar _gv_i_154;
											for (_gv_i_154 = 0; _gv_i_154 < NUM_LANES; _gv_i_154 = _gv_i_154 + 1) begin : g_rs1_data
												localparam i = _gv_i_154;
												// Trace: src/VX_csr_unit.sv:33:9
												assign rs1_data[i * 32+:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[259 + (i * 32)+:32];
											end
											// Trace: src/VX_csr_unit.sv:35:5
											localparam VX_gpu_pkg_INST_SFU_CSRRW = 4'h6;
											wire csr_write_enable = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[433-:4] == VX_gpu_pkg_INST_SFU_CSRRW;
											// Trace: src/VX_csr_unit.sv:36:5
											// expanded module instance: csr_data
											localparam _param_9D0B6_INSTANCE_ID = INSTANCE_ID;
											localparam _param_9D0B6_CORE_ID = CORE_ID;
											if (1) begin : csr_data
												// removed import VX_gpu_pkg::*;
												// Trace: src/VX_csr_data.sv:4:15
												localparam INSTANCE_ID = _param_9D0B6_INSTANCE_ID;
												// Trace: src/VX_csr_data.sv:5:15
												localparam CORE_ID = _param_9D0B6_CORE_ID;
												// Trace: src/VX_csr_data.sv:7:5
												wire clk;
												// Trace: src/VX_csr_data.sv:8:5
												wire reset;
												// Trace: src/VX_csr_data.sv:9:5
												// removed localparam type VX_gpu_pkg_base_dcrs_t
												wire [71:0] base_dcrs;
												// Trace: src/VX_csr_data.sv:10:5
												// removed modport instance commit_csr_if
												// Trace: src/VX_csr_data.sv:11:5
												localparam VX_gpu_pkg_PERF_CTR_BITS = 44;
												wire [43:0] cycles;
												// Trace: src/VX_csr_data.sv:12:5
												wire [3:0] active_warps;
												// Trace: src/VX_csr_data.sv:13:5
												wire [15:0] thread_masks;
												// Trace: src/VX_csr_data.sv:14:5
												wire read_enable;
												// Trace: src/VX_csr_data.sv:15:5
												localparam VX_gpu_pkg_UUID_WIDTH = 1;
												wire [0:0] read_uuid;
												// Trace: src/VX_csr_data.sv:16:5
												localparam VX_gpu_pkg_NW_BITS = 2;
												localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
												wire [1:0] read_wid;
												// Trace: src/VX_csr_data.sv:17:5
												wire [11:0] read_addr;
												// Trace: src/VX_csr_data.sv:18:5
												wire [31:0] read_data_ro;
												// Trace: src/VX_csr_data.sv:19:5
												wire [31:0] read_data_rw;
												// Trace: src/VX_csr_data.sv:20:5
												wire write_enable;
												// Trace: src/VX_csr_data.sv:21:5
												wire [0:0] write_uuid;
												// Trace: src/VX_csr_data.sv:22:5
												wire [1:0] write_wid;
												// Trace: src/VX_csr_data.sv:23:5
												wire [11:0] write_addr;
												// Trace: src/VX_csr_data.sv:24:5
												wire [31:0] write_data;
												// Trace: src/VX_csr_data.sv:26:5
												reg [31:0] mscratch;
												// Trace: src/VX_csr_data.sv:27:5
												always @(posedge clk) begin
													// Trace: src/VX_csr_data.sv:28:9
													if (reset)
														// Trace: src/VX_csr_data.sv:29:13
														mscratch <= base_dcrs[39-:32];
													if (write_enable)
														// Trace: src/VX_csr_data.sv:32:13
														case (write_addr)
															12'h180, 12'h300, 12'h744, 12'h302, 12'h303, 12'h304, 12'h305, 12'h341, 12'h3a0, 12'h3b0:
																;
															12'h340:
																// Trace: src/VX_csr_data.sv:45:21
																mscratch <= write_data;
															default:
																;
														endcase
												end
												// Trace: src/VX_csr_data.sv:53:5
												reg [31:0] read_data_ro_w;
												// Trace: src/VX_csr_data.sv:54:5
												reg [31:0] read_data_rw_w;
												// Trace: src/VX_csr_data.sv:55:5
												reg read_addr_valid_w;
												// Trace: src/VX_csr_data.sv:56:5
												always @(*) begin
													// Trace: src/VX_csr_data.sv:57:9
													read_data_ro_w = 1'sb0;
													// Trace: src/VX_csr_data.sv:58:9
													read_data_rw_w = 1'sb0;
													// Trace: src/VX_csr_data.sv:59:9
													read_addr_valid_w = 1;
													// Trace: src/VX_csr_data.sv:60:9
													case (read_addr)
														12'hf11:
															// Trace: src/VX_csr_data.sv:61:24
															read_data_ro_w = 32'sd0;
														12'hf12:
															// Trace: src/VX_csr_data.sv:62:26
															read_data_ro_w = 32'sd0;
														12'hf13:
															// Trace: src/VX_csr_data.sv:63:27
															read_data_ro_w = 32'sd0;
														12'h301:
															// Trace: src/VX_csr_data.sv:64:29
															read_data_ro_w = 32'h40901100;
														12'h340:
															// Trace: src/VX_csr_data.sv:90:25
															read_data_rw_w = mscratch;
														12'hcc1:
															// Trace: src/VX_csr_data.sv:91:26
															read_data_ro_w = sv2v_cast_32(read_wid);
														12'hcc2:
															// Trace: src/VX_csr_data.sv:92:26
															read_data_ro_w = sv2v_cast_32_signed(CORE_ID);
														12'hcc4:
															// Trace: src/VX_csr_data.sv:93:22
															read_data_ro_w = sv2v_cast_32(thread_masks[read_wid * 4+:4]);
														12'hcc3:
															// Trace: src/VX_csr_data.sv:94:22
															read_data_ro_w = sv2v_cast_32(active_warps);
														12'hfc0:
															// Trace: src/VX_csr_data.sv:95:22
															read_data_ro_w = 32'sd4;
														12'hfc1:
															// Trace: src/VX_csr_data.sv:96:24
															read_data_ro_w = 32'sd4;
														12'hfc2:
															// Trace: src/VX_csr_data.sv:97:24
															read_data_ro_w = 32'sd1;
														12'hfc3:
															// Trace: src/VX_csr_data.sv:98:22
															read_data_ro_w = 32'hffff0000;
														12'hb00:
															// Trace: src/VX_csr_data.sv:99:19
															read_data_ro_w = cycles[31:0];
														12'hb00 + 12'h080:
															// Trace: src/VX_csr_data.sv:100:26
															read_data_ro_w = sv2v_cast_32(cycles[43:32]);
														12'hb01:
															// Trace: src/VX_csr_data.sv:101:23
															read_data_ro_w = 1'sbx;
														12'hb81:
															// Trace: src/VX_csr_data.sv:102:23
															read_data_ro_w = 1'sbx;
														12'hb02:
															// Trace: src/VX_csr_data.sv:103:19
															read_data_ro_w = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_csr_if.instret[31:0];
														12'hb02 + 12'h080:
															// Trace: src/VX_csr_data.sv:104:26
															read_data_ro_w = sv2v_cast_32(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_csr_if.instret[43:32]);
														12'h180, 12'h300, 12'h744, 12'h302, 12'h303, 12'h304, 12'h305, 12'h341, 12'h3a0, 12'h3b0:
															// Trace: src/VX_csr_data.sv:114:23
															read_data_ro_w = 32'sd0;
														default: begin
															// Trace: src/VX_csr_data.sv:116:17
															read_addr_valid_w = 0;
															// Trace: src/VX_csr_data.sv:117:17
															if (((read_addr >= 12'hb03) && (read_addr < 2851)) || ((read_addr >= 12'hb83) && (read_addr < 2979)))
																// Trace: src/VX_csr_data.sv:119:21
																read_addr_valid_w = 1;
														end
													endcase
												end
												// Trace: src/VX_csr_data.sv:124:5
												assign read_data_ro = read_data_ro_w;
												// Trace: src/VX_csr_data.sv:125:5
												assign read_data_rw = read_data_rw_w;
											end
											assign csr_data.clk = clk;
											assign csr_data.reset = reset;
											assign csr_data.base_dcrs = base_dcrs;
											assign csr_data.cycles = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.cycles;
											assign csr_data.active_warps = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.active_warps;
											assign csr_data.thread_masks = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.thread_masks;
											assign csr_data.read_enable = csr_req_valid && csr_rd_enable;
											assign csr_data.read_uuid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[470];
											assign csr_data.read_wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[469-:2];
											assign csr_data.read_addr = csr_addr;
											assign csr_read_data_ro = csr_data.read_data_ro;
											assign csr_read_data_rw = csr_data.read_data_rw;
											assign csr_data.write_enable = csr_req_valid && csr_wr_enable;
											assign csr_data.write_uuid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[470];
											assign csr_data.write_wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[469-:2];
											assign csr_data.write_addr = csr_addr;
											assign csr_data.write_data = csr_write_data;
											// Trace: src/VX_csr_unit.sv:59:5
											wire [127:0] wtid;
											wire [127:0] gtid;
											// Trace: src/VX_csr_unit.sv:60:5
											genvar _gv_i_155;
											for (_gv_i_155 = 0; _gv_i_155 < NUM_LANES; _gv_i_155 = _gv_i_155 + 1) begin : g_wtid
												localparam i = _gv_i_155;
												if (1) begin : g_no_pid
													// Trace: src/VX_csr_unit.sv:64:13
													assign wtid[i * 32+:32] = i;
												end
											end
											// Trace: src/VX_csr_unit.sv:67:5
											genvar _gv_i_156;
											localparam VX_gpu_pkg_NT_BITS = 2;
											for (_gv_i_156 = 0; _gv_i_156 < NUM_LANES; _gv_i_156 = _gv_i_156 + 1) begin : g_gtid
												localparam i = _gv_i_156;
												// Trace: src/VX_csr_unit.sv:68:9
												assign gtid[i * 32+:32] = ((sv2v_cast_32_signed(CORE_ID) << 4) + (sv2v_cast_32(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[469-:2]) << VX_gpu_pkg_NT_BITS)) + wtid[i * 32+:32];
											end
											// Trace: src/VX_csr_unit.sv:70:5
											always @(*) begin
												// Trace: src/VX_csr_unit.sv:71:9
												csr_rd_enable = 0;
												// Trace: src/VX_csr_unit.sv:72:9
												case (csr_addr)
													12'hcc0:
														// Trace: src/VX_csr_unit.sv:73:19
														csr_read_data = wtid;
													12'hf14:
														// Trace: src/VX_csr_unit.sv:74:21
														csr_read_data = gtid;
													default: begin
														// Trace: src/VX_csr_unit.sv:76:13
														csr_read_data = {NUM_LANES {csr_read_data_ro | csr_read_data_rw}};
														// Trace: src/VX_csr_unit.sv:77:13
														csr_rd_enable = 1;
													end
												endcase
											end
											// Trace: src/VX_csr_unit.sv:81:5
											assign csr_req_data = (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[410] ? sv2v_cast_32(csr_imm) : rs1_data[0+:32]);
											// Trace: src/VX_csr_unit.sv:82:5
											assign csr_wr_enable = csr_write_enable || |csr_req_data;
											// Trace: src/VX_csr_unit.sv:83:5
											localparam VX_gpu_pkg_INST_SFU_CSRRS = 4'h7;
											always @(*)
												// Trace: src/VX_csr_unit.sv:84:9
												case (Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[433-:4])
													VX_gpu_pkg_INST_SFU_CSRRW:
														// Trace: src/VX_csr_unit.sv:86:17
														csr_write_data = csr_req_data;
													VX_gpu_pkg_INST_SFU_CSRRS:
														// Trace: src/VX_csr_unit.sv:89:17
														csr_write_data = csr_read_data_rw | csr_req_data;
													default:
														// Trace: src/VX_csr_unit.sv:92:17
														csr_write_data = csr_read_data_rw & ~csr_req_data;
												endcase
											// Trace: src/VX_csr_unit.sv:96:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.unlock_warp = ((csr_req_valid && csr_req_ready) && Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[0]) && is_fpu_csr;
											// Trace: src/VX_csr_unit.sv:97:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.sched_csr_if.unlock_wid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[469-:2];
											// Trace: src/VX_csr_unit.sv:98:5
											VX_elastic_buffer #(
												.DATAW(DATAW),
												.SIZE(2)
											) rsp_buf(
												.clk(clk),
												.reset(reset),
												.valid_in(csr_req_valid),
												.ready_in(csr_req_ready),
												.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[470], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[469-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[467-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[463-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[391-:5], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[392], csr_read_data, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_execute_if[_mbase_execute_if].data[0]}),
												.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[173], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[172-:2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[170-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[166-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[135-:5], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[136], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[130-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[2], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[1], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].data[0]}),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].valid),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.pe_result_if[_mbase_result_if].ready)
											);
										end
										assign csr_unit.clk = clk;
										assign csr_unit.reset = reset;
										assign csr_unit.base_dcrs = base_dcrs;
										// Trace: src/VX_sfu_unit.sv:87:5
										// expanded module instance: gather_unit
										localparam _bbase_8E516_result_if = 0;
										localparam _bbase_8E516_commit_if = 2;
										localparam _param_8E516_BLOCK_SIZE = BLOCK_SIZE;
										localparam _param_8E516_NUM_LANES = NUM_LANES;
										localparam _param_8E516_OUT_BUF = 3;
										if (1) begin : gather_unit
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_gather_unit.sv:2:15
											localparam BLOCK_SIZE = _param_8E516_BLOCK_SIZE;
											// Trace: src/VX_gather_unit.sv:3:15
											localparam NUM_LANES = _param_8E516_NUM_LANES;
											// Trace: src/VX_gather_unit.sv:4:15
											localparam OUT_BUF = _param_8E516_OUT_BUF;
											// Trace: src/VX_gather_unit.sv:6:5
											wire clk;
											// Trace: src/VX_gather_unit.sv:7:5
											wire reset;
											// Trace: src/VX_gather_unit.sv:8:5
											localparam _mbase_result_if = 0;
											// Trace: src/VX_gather_unit.sv:9:5
											localparam _mbase_commit_if = 2;
											// Trace: src/VX_gather_unit.sv:11:5
											localparam BLOCK_SIZE_W = 1;
											// Trace: src/VX_gather_unit.sv:12:5
											localparam NUM_PACKETS = 1;
											// Trace: src/VX_gather_unit.sv:13:5
											localparam LPID_BITS = 0;
											// Trace: src/VX_gather_unit.sv:14:5
											localparam LPID_WIDTH = 1;
											// Trace: src/VX_gather_unit.sv:15:5
											localparam GPID_BITS = 0;
											// Trace: src/VX_gather_unit.sv:16:5
											localparam GPID_WIDTH = 1;
											// Trace: src/VX_gather_unit.sv:17:5
											localparam VX_gpu_pkg_REG_TYPES = 1;
											localparam VX_gpu_pkg_RV_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS = 32;
											localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
											localparam VX_gpu_pkg_NW_BITS = 2;
											localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
											localparam VX_gpu_pkg_PC_BITS = 30;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam DATAW = 174;
											// Trace: src/VX_gather_unit.sv:18:5
											localparam DATA_WIS_OFF = 171;
											// Trace: src/VX_gather_unit.sv:19:5
											wire [0:0] result_in_valid;
											// Trace: src/VX_gather_unit.sv:20:5
											wire [173:0] result_in_data;
											// Trace: src/VX_gather_unit.sv:21:5
											wire [0:0] result_in_ready;
											// Trace: src/VX_gather_unit.sv:22:5
											localparam VX_gpu_pkg_ISSUE_ISW_BITS = 0;
											localparam VX_gpu_pkg_ISSUE_ISW_W = 1;
											wire [0:0] result_in_isw;
											// Trace: src/VX_gather_unit.sv:23:5
											genvar _gv_i_60;
											for (_gv_i_60 = 0; _gv_i_60 < BLOCK_SIZE; _gv_i_60 = _gv_i_60 + 1) begin : g_commit_in
												localparam i = _gv_i_60;
												// Trace: src/VX_gather_unit.sv:24:9
												assign result_in_valid[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_result_if[i + _mbase_result_if].valid;
												// Trace: src/VX_gather_unit.sv:25:9
												assign result_in_data[i * 174+:174] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_result_if[i + _mbase_result_if].data;
												// Trace: src/VX_gather_unit.sv:26:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.execute.sfu_unit.per_block_result_if[i + _mbase_result_if].ready = result_in_ready[i];
												if (1) begin : g_result_in_isw_full
													// Trace: src/VX_gather_unit.sv:34:13
													assign result_in_isw[i+:1] = sv2v_cast_1_signed(i);
												end
											end
											// Trace: src/VX_gather_unit.sv:37:5
											reg [0:0] result_out_valid;
											// Trace: src/VX_gather_unit.sv:38:5
											reg [173:0] result_out_data;
											// Trace: src/VX_gather_unit.sv:39:5
											wire [0:0] result_out_ready;
											// Trace: src/VX_gather_unit.sv:40:5
											always @(*) begin
												// Trace: src/VX_gather_unit.sv:41:9
												result_out_valid = 1'sb0;
												// Trace: src/VX_gather_unit.sv:42:9
												begin : sv2v_autoblock_15
													// Trace: src/VX_gather_unit.sv:42:14
													integer i;
													// Trace: src/VX_gather_unit.sv:42:14
													for (i = 0; i < 1; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:43:13
															result_out_data[i * 174+:174] = 1'sbx;
														end
												end
												begin : sv2v_autoblock_16
													// Trace: src/VX_gather_unit.sv:45:14
													integer i;
													// Trace: src/VX_gather_unit.sv:45:14
													for (i = 0; i < BLOCK_SIZE; i = i + 1)
														begin
															// Trace: src/VX_gather_unit.sv:46:13
															result_out_valid[result_in_isw[i+:1]] = result_in_valid[i];
															// Trace: src/VX_gather_unit.sv:47:13
															result_out_data[result_in_isw[i+:1] * 174+:174] = result_in_data[i * 174+:174];
														end
												end
											end
											// Trace: src/VX_gather_unit.sv:50:5
											genvar _gv_i_61;
											for (_gv_i_61 = 0; _gv_i_61 < BLOCK_SIZE; _gv_i_61 = _gv_i_61 + 1) begin : g_result_in_ready
												localparam i = _gv_i_61;
												// Trace: src/VX_gather_unit.sv:51:9
												assign result_in_ready[i] = result_out_ready[result_in_isw[i+:1]];
											end
											// Trace: src/VX_gather_unit.sv:53:5
											genvar _gv_i_62;
											localparam VX_gpu_pkg_SIMD_COUNT = 1;
											localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
											localparam VX_gpu_pkg_SIMD_IDX_W = 1;
											for (_gv_i_62 = 0; _gv_i_62 < 1; _gv_i_62 = _gv_i_62 + 1) begin : g_out_bufs
												localparam i = _gv_i_62;
												// Trace: src/VX_gather_unit.sv:54:9
												// expanded interface instance: result_tmp_if
												localparam _param_D4A7C_NUM_LANES = NUM_LANES;
												if (1) begin : result_tmp_if
													// removed import VX_gpu_pkg::*;
													// Trace: src/VX_result_if.sv:2:15
													localparam NUM_LANES = _param_D4A7C_NUM_LANES;
													// Trace: src/VX_result_if.sv:3:15
													localparam PID_WIDTH = 1;
													// Trace: src/VX_result_if.sv:5:5
													localparam VX_gpu_pkg_REG_TYPES = 1;
													localparam VX_gpu_pkg_RV_REGS = 32;
													localparam VX_gpu_pkg_NUM_REGS = 32;
													localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
													localparam VX_gpu_pkg_NW_BITS = 2;
													localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
													localparam VX_gpu_pkg_PC_BITS = 30;
													localparam VX_gpu_pkg_UUID_WIDTH = 1;
													// removed localparam type data_t
													// Trace: src/VX_result_if.sv:17:5
													wire valid;
													// Trace: src/VX_result_if.sv:18:5
													wire [173:0] data;
													// Trace: src/VX_result_if.sv:19:5
													wire ready;
													// Trace: src/VX_result_if.sv:20:5
													// Trace: src/VX_result_if.sv:25:5
												end
												// Trace: src/VX_gather_unit.sv:57:9
												VX_elastic_buffer #(
													.DATAW(DATAW),
													.SIZE(2),
													.OUT_REG(1)
												) out_buf(
													.clk(clk),
													.reset(reset),
													.valid_in(result_out_valid[i]),
													.ready_in(result_out_ready[i]),
													.data_in(result_out_data[i * 174+:174]),
													.data_out(result_tmp_if.data),
													.valid_out(result_tmp_if.valid),
													.ready_out(result_tmp_if.ready)
												);
												// Trace: src/VX_gather_unit.sv:71:9
												wire [0:0] commit_sid_w;
												// Trace: src/VX_gather_unit.sv:72:9
												wire [3:0] commit_tmask_w;
												// Trace: src/VX_gather_unit.sv:73:9
												wire [127:0] commit_data_w;
												if (1) begin : g_no_lpid
													// Trace: src/VX_gather_unit.sv:91:13
													assign commit_sid_w = result_tmp_if.data[2];
													// Trace: src/VX_gather_unit.sv:92:13
													assign commit_tmask_w = result_tmp_if.data[170-:4];
													// Trace: src/VX_gather_unit.sv:93:13
													assign commit_data_w = result_tmp_if.data[130-:128];
												end
												// Trace: src/VX_gather_unit.sv:95:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_if].valid = result_tmp_if.valid;
												// Trace: src/VX_gather_unit.sv:96:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_if].data = {result_tmp_if.data[173], result_tmp_if.data[172-:2], commit_sid_w, commit_tmask_w, result_tmp_if.data[166-:30], result_tmp_if.data[136], result_tmp_if.data[135-:5], commit_data_w, result_tmp_if.data[1], result_tmp_if.data[0]};
												// Trace: src/VX_gather_unit.sv:108:9
												assign result_tmp_if.ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[i + _mbase_commit_if].ready;
											end
										end
										assign gather_unit.clk = clk;
										assign gather_unit.reset = reset;
									end
									assign sfu_unit.clk = clk;
									assign sfu_unit.reset = reset;
									assign sfu_unit.base_dcrs = base_dcrs;
								end
								assign execute.clk = clk;
								assign execute.reset = reset;
								assign execute.base_dcrs = base_dcrs;
								// Trace: src/VX_core.sv:97:5
								// expanded module instance: commit
								localparam _bbase_D837E_commit_if = 0;
								localparam _bbase_D837E_writeback_if = 0;
								localparam _param_D837E_INSTANCE_ID = "";
								if (1) begin : commit
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_commit.sv:2:15
									localparam INSTANCE_ID = _param_D837E_INSTANCE_ID;
									// Trace: src/VX_commit.sv:4:5
									wire clk;
									// Trace: src/VX_commit.sv:5:5
									wire reset;
									// Trace: src/VX_commit.sv:6:5
									localparam VX_gpu_pkg_EX_SFU = 2;
									localparam VX_gpu_pkg_EX_FPU = 2;
									localparam VX_gpu_pkg_EX_TCU = 2;
									localparam VX_gpu_pkg_NUM_EX_UNITS = 3;
									localparam _mbase_commit_if = 0;
									// Trace: src/VX_commit.sv:7:5
									localparam _mbase_writeback_if = 0;
									// Trace: src/VX_commit.sv:8:5
									// removed modport instance commit_csr_if
									// Trace: src/VX_commit.sv:9:5
									// removed modport instance commit_sched_if
									// Trace: src/VX_commit.sv:11:5
									localparam VX_gpu_pkg_REG_TYPES = 1;
									localparam VX_gpu_pkg_RV_REGS = 32;
									localparam VX_gpu_pkg_NUM_REGS = 32;
									localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
									localparam VX_gpu_pkg_NW_BITS = 2;
									localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
									localparam VX_gpu_pkg_PC_BITS = 30;
									localparam VX_gpu_pkg_SIMD_COUNT = 1;
									localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
									localparam VX_gpu_pkg_SIMD_IDX_W = 1;
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									// removed localparam type VX_gpu_pkg_commit_t
									localparam OUT_DATAW = 174;
									// Trace: src/VX_commit.sv:12:5
									localparam COMMIT_SIZEW = 3;
									// Trace: src/VX_commit.sv:13:5
									localparam COMMIT_ALL_SIZEW = 3;
									// Trace: src/VX_commit.sv:14:5
									// expanded interface instance: commit_arb_if
									genvar _arr_25972;
									for (_arr_25972 = 0; _arr_25972 <= 0; _arr_25972 = _arr_25972 + 1) begin : commit_arb_if
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_commit_if.sv:2:5
										wire valid;
										// Trace: src/VX_commit_if.sv:3:5
										localparam VX_gpu_pkg_REG_TYPES = 1;
										localparam VX_gpu_pkg_RV_REGS = 32;
										localparam VX_gpu_pkg_NUM_REGS = 32;
										localparam VX_gpu_pkg_NUM_REGS_BITS = 5;
										localparam VX_gpu_pkg_NW_BITS = 2;
										localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
										localparam VX_gpu_pkg_PC_BITS = 30;
										localparam VX_gpu_pkg_SIMD_COUNT = 1;
										localparam VX_gpu_pkg_SIMD_IDX_BITS = 0;
										localparam VX_gpu_pkg_SIMD_IDX_W = 1;
										localparam VX_gpu_pkg_UUID_WIDTH = 1;
										// removed localparam type VX_gpu_pkg_commit_t
										wire [173:0] data;
										// Trace: src/VX_commit_if.sv:4:5
										wire ready;
										// Trace: src/VX_commit_if.sv:5:5
										// Trace: src/VX_commit_if.sv:10:5
									end
									// Trace: src/VX_commit.sv:15:5
									wire [0:0] per_issue_commit_fire;
									// Trace: src/VX_commit.sv:16:5
									wire [1:0] per_issue_commit_wid;
									// Trace: src/VX_commit.sv:17:5
									wire [3:0] per_issue_commit_tmask;
									// Trace: src/VX_commit.sv:18:5
									wire [0:0] per_issue_commit_eop;
									// Trace: src/VX_commit.sv:19:5
									genvar _gv_i_80;
									for (_gv_i_80 = 0; _gv_i_80 < 1; _gv_i_80 = _gv_i_80 + 1) begin : g_commit_arbs
										localparam i = _gv_i_80;
										// Trace: src/VX_commit.sv:20:9
										wire [2:0] valid_in;
										// Trace: src/VX_commit.sv:21:9
										wire [521:0] data_in;
										// Trace: src/VX_commit.sv:22:9
										wire [2:0] ready_in;
										genvar _gv_j_12;
										for (_gv_j_12 = 0; _gv_j_12 < VX_gpu_pkg_NUM_EX_UNITS; _gv_j_12 = _gv_j_12 + 1) begin : g_data_in
											localparam j = _gv_j_12;
											// Trace: src/VX_commit.sv:24:13
											assign valid_in[j] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[((j * 1) + i) + _mbase_commit_if].valid;
											// Trace: src/VX_commit.sv:25:13
											assign data_in[j * 174+:174] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[((j * 1) + i) + _mbase_commit_if].data;
											// Trace: src/VX_commit.sv:26:13
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_if[((j * 1) + i) + _mbase_commit_if].ready = ready_in[j];
										end
										// Trace: src/VX_commit.sv:28:9
										VX_stream_arb #(
											.NUM_INPUTS(VX_gpu_pkg_NUM_EX_UNITS),
											.DATAW(OUT_DATAW),
											.ARBITER("P"),
											.OUT_BUF(1)
										) commit_arb(
											.clk(clk),
											.reset(reset),
											.valid_in(valid_in),
											.ready_in(ready_in),
											.data_in(data_in),
											.data_out(commit_arb_if[i].data),
											.valid_out(commit_arb_if[i].valid),
											.ready_out(commit_arb_if[i].ready),
											.sel_out()
										);
										// Trace: src/VX_commit.sv:44:9
										assign per_issue_commit_fire[i] = commit_arb_if[i].valid && commit_arb_if[i].ready;
										// Trace: src/VX_commit.sv:45:9
										assign per_issue_commit_tmask[i * 4+:4] = {4 {per_issue_commit_fire[i]}} & commit_arb_if[i].data[169-:4];
										// Trace: src/VX_commit.sv:46:9
										assign per_issue_commit_wid[i * 2+:2] = commit_arb_if[i].data[172-:2];
										// Trace: src/VX_commit.sv:47:9
										assign per_issue_commit_eop[i] = commit_arb_if[i].data[0];
									end
									// Trace: src/VX_commit.sv:49:5
									wire [2:0] commit_size;
									wire [2:0] commit_size_r;
									// Trace: src/VX_commit.sv:50:5
									wire [2:0] commit_size_all_r;
									wire [2:0] commit_size_all_rr;
									// Trace: src/VX_commit.sv:51:5
									wire commit_fire_any;
									wire commit_fire_any_r;
									wire commit_fire_any_rr;
									// Trace: src/VX_commit.sv:52:5
									assign commit_fire_any = |per_issue_commit_fire;
									// Trace: src/VX_commit.sv:53:5
									genvar _gv_i_81;
									for (_gv_i_81 = 0; _gv_i_81 < 1; _gv_i_81 = _gv_i_81 + 1) begin : g_commit_size
										localparam i = _gv_i_81;
										// Trace: src/VX_commit.sv:54:9
										wire [2:0] count;
										// Trace: src/VX_commit.sv:55:5
										VX_popcount #(
											.N(4),
											.MODEL(1)
										) __pop_count_ex89(
											.data_in(per_issue_commit_tmask[i * 4+:4]),
											.data_out(count)
										);
										// Trace: src/VX_commit.sv:62:9
										assign commit_size[i * 3+:3] = count;
									end
									// Trace: src/VX_commit.sv:64:5
									VX_pipe_register #(
										.DATAW(4),
										.RESETW(1)
									) commit_size_reg1(
										.clk(clk),
										.reset(reset),
										.enable(1'b1),
										.data_in({commit_fire_any, commit_size}),
										.data_out({commit_fire_any_r, commit_size_r})
									);
									// Trace: src/VX_commit.sv:74:5
									VX_reduce_tree #(
										.DATAW_IN(COMMIT_SIZEW),
										.DATAW_OUT(COMMIT_ALL_SIZEW),
										.N(1),
										.OP("+")
									) commit_size_reduce(
										.data_in(commit_size_r),
										.data_out(commit_size_all_r)
									);
									// Trace: src/VX_commit.sv:83:5
									VX_pipe_register #(
										.DATAW(4),
										.RESETW(1)
									) commit_size_reg2(
										.clk(clk),
										.reset(reset),
										.enable(1'b1),
										.data_in({commit_fire_any_r, commit_size_all_r}),
										.data_out({commit_fire_any_rr, commit_size_all_rr})
									);
									// Trace: src/VX_commit.sv:93:5
									localparam VX_gpu_pkg_PERF_CTR_BITS = 44;
									reg [43:0] instret;
									// Trace: src/VX_commit.sv:94:5
									always @(posedge clk)
										// Trace: src/VX_commit.sv:95:8
										if (reset)
											// Trace: src/VX_commit.sv:96:13
											instret <= 1'sb0;
										else
											// Trace: src/VX_commit.sv:98:13
											if (commit_fire_any_rr)
												// Trace: src/VX_commit.sv:99:17
												instret <= instret + sv2v_cast_44(commit_size_all_rr);
									// Trace: src/VX_commit.sv:103:5
									assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_csr_if.instret = instret;
									// Trace: src/VX_commit.sv:104:5
									reg [3:0] committed_warps;
									// Trace: src/VX_commit.sv:105:5
									always @(*) begin
										// Trace: src/VX_commit.sv:106:9
										committed_warps = 0;
										// Trace: src/VX_commit.sv:107:9
										begin : sv2v_autoblock_17
											// Trace: src/VX_commit.sv:107:14
											integer i;
											// Trace: src/VX_commit.sv:107:14
											for (i = 0; i < 1; i = i + 1)
												begin
													// Trace: src/VX_commit.sv:108:13
													if (per_issue_commit_fire[i] && per_issue_commit_eop[i])
														// Trace: src/VX_commit.sv:109:17
														committed_warps[per_issue_commit_wid[i * 2+:2]] = 1;
												end
										end
									end
									// Trace: src/VX_commit.sv:113:5
									VX_pipe_register #(
										.DATAW(4),
										.RESETW(4)
									) committed_pipe_reg(
										.clk(clk),
										.reset(reset),
										.enable(1'b1),
										.data_in(committed_warps),
										.data_out({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.commit_sched_if.committed_warps})
									);
									// Trace: src/VX_commit.sv:123:5
									genvar _gv_i_82;
									localparam VX_gpu_pkg_ISSUE_ISW_BITS = 0;
									localparam VX_gpu_pkg_PER_ISSUE_WARPS = 4;
									localparam VX_gpu_pkg_ISSUE_WIS_BITS = 2;
									localparam VX_gpu_pkg_ISSUE_WIS_W = VX_gpu_pkg_ISSUE_WIS_BITS;
									function automatic [1:0] VX_gpu_pkg_wid_to_wis;
										// Trace: src/VX_gpu_pkg.sv:285:9
										input reg [1:0] wid;
										// Trace: src/VX_gpu_pkg.sv:287:9
										begin
											// Trace: src/VX_gpu_pkg.sv:288:13
											VX_gpu_pkg_wid_to_wis = wid >> VX_gpu_pkg_ISSUE_ISW_BITS;
										end
									endfunction
									for (_gv_i_82 = 0; _gv_i_82 < 1; _gv_i_82 = _gv_i_82 + 1) begin : g_writeback
										localparam i = _gv_i_82;
										// Trace: src/VX_commit.sv:124:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].valid = commit_arb_if[i].valid && commit_arb_if[i].data[135];
										// Trace: src/VX_commit.sv:125:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[172] = commit_arb_if[i].data[173];
										// Trace: src/VX_commit.sv:126:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[171-:2] = VX_gpu_pkg_wid_to_wis(commit_arb_if[i].data[172-:2]);
										// Trace: src/VX_commit.sv:127:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[169] = commit_arb_if[i].data[170];
										// Trace: src/VX_commit.sv:128:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[164-:30] = commit_arb_if[i].data[165-:30];
										// Trace: src/VX_commit.sv:129:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[168-:4] = commit_arb_if[i].data[169-:4];
										// Trace: src/VX_commit.sv:130:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[134-:5] = commit_arb_if[i].data[134-:5];
										// Trace: src/VX_commit.sv:131:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[129-:128] = commit_arb_if[i].data[129-:128];
										// Trace: src/VX_commit.sv:132:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[1] = commit_arb_if[i].data[1];
										// Trace: src/VX_commit.sv:133:9
										assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.writeback_if[i + _mbase_writeback_if].data[0] = commit_arb_if[i].data[0];
										// Trace: src/VX_commit.sv:134:9
										assign commit_arb_if[i].ready = 1;
									end
								end
								assign commit.clk = clk;
								assign commit.reset = reset;
								// Trace: src/VX_core.sv:107:5
								// expanded module instance: mem_unit
								localparam _bbase_A06D0_lsu_mem_if = 0;
								localparam _bbase_A06D0_dcache_bus_if = core_id * VX_gpu_pkg_DCACHE_NUM_REQS;
								localparam _param_A06D0_INSTANCE_ID = INSTANCE_ID;
								if (1) begin : mem_unit
									// removed import VX_gpu_pkg::*;
									// Trace: src/VX_mem_unit.sv:2:15
									localparam INSTANCE_ID = _param_A06D0_INSTANCE_ID;
									// Trace: src/VX_mem_unit.sv:4:5
									wire clk;
									// Trace: src/VX_mem_unit.sv:5:5
									wire reset;
									// Trace: src/VX_mem_unit.sv:6:5
									localparam _mbase_lsu_mem_if = 0;
									// Trace: src/VX_mem_unit.sv:7:5
									localparam VX_gpu_pkg_DCACHE_WORD_SIZE = 16;
									localparam VX_gpu_pkg_XLENB = 4;
									localparam VX_gpu_pkg_LSU_WORD_SIZE = VX_gpu_pkg_XLENB;
									localparam VX_gpu_pkg_DCACHE_CHANNELS = 1;
									localparam VX_gpu_pkg_DCACHE_NUM_REQS = 1;
									localparam _mbase_dcache_bus_if = _bbase_A06D0_dcache_bus_if;
									// Trace: src/VX_mem_unit.sv:9:5
									localparam VX_gpu_pkg_LSU_MEM_BATCHES = 1;
									localparam VX_gpu_pkg_LSU_TAG_ID_BITS = 1;
									localparam VX_gpu_pkg_UUID_WIDTH = 1;
									localparam VX_gpu_pkg_LSU_TAG_WIDTH = 2;
									// expanded interface instance: lsu_dcache_if
									localparam _param_9E566_NUM_LANES = 4;
									localparam _param_9E566_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
									localparam _param_9E566_TAG_WIDTH = VX_gpu_pkg_LSU_TAG_WIDTH;
									genvar _arr_9E566;
									for (_arr_9E566 = 0; _arr_9E566 <= 0; _arr_9E566 = _arr_9E566 + 1) begin : lsu_dcache_if
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_lsu_mem_if.sv:2:15
										localparam NUM_LANES = _param_9E566_NUM_LANES;
										// Trace: src/VX_lsu_mem_if.sv:3:15
										localparam DATA_SIZE = _param_9E566_DATA_SIZE;
										// Trace: src/VX_lsu_mem_if.sv:4:15
										localparam TAG_WIDTH = _param_9E566_TAG_WIDTH;
										// Trace: src/VX_lsu_mem_if.sv:5:15
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
										// Trace: src/VX_lsu_mem_if.sv:6:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_lsu_mem_if.sv:7:15
										localparam ADDR_WIDTH = 30;
										// Trace: src/VX_lsu_mem_if.sv:9:5
										localparam VX_gpu_pkg_UUID_WIDTH = 1;
										// removed localparam type tag_t
										// Trace: src/VX_lsu_mem_if.sv:13:5
										// removed localparam type req_data_t
										// Trace: src/VX_lsu_mem_if.sv:22:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_lsu_mem_if.sv:27:5
										wire req_valid;
										// Trace: src/VX_lsu_mem_if.sv:28:5
										wire [282:0] req_data;
										// Trace: src/VX_lsu_mem_if.sv:29:5
										wire req_ready;
										// Trace: src/VX_lsu_mem_if.sv:30:5
										wire rsp_valid;
										// Trace: src/VX_lsu_mem_if.sv:31:5
										wire [133:0] rsp_data;
										// Trace: src/VX_lsu_mem_if.sv:32:5
										wire rsp_ready;
										// Trace: src/VX_lsu_mem_if.sv:33:5
										// Trace: src/VX_lsu_mem_if.sv:41:5
									end
									// Trace: src/VX_mem_unit.sv:14:5
									localparam LMEM_ADDR_WIDTH = 12;
									// Trace: src/VX_mem_unit.sv:15:5
									// expanded interface instance: lsu_lmem_if
									localparam _param_B7A65_NUM_LANES = 4;
									localparam _param_B7A65_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
									localparam _param_B7A65_TAG_WIDTH = VX_gpu_pkg_LSU_TAG_WIDTH;
									genvar _arr_B7A65;
									for (_arr_B7A65 = 0; _arr_B7A65 <= 0; _arr_B7A65 = _arr_B7A65 + 1) begin : lsu_lmem_if
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_lsu_mem_if.sv:2:15
										localparam NUM_LANES = _param_B7A65_NUM_LANES;
										// Trace: src/VX_lsu_mem_if.sv:3:15
										localparam DATA_SIZE = _param_B7A65_DATA_SIZE;
										// Trace: src/VX_lsu_mem_if.sv:4:15
										localparam TAG_WIDTH = _param_B7A65_TAG_WIDTH;
										// Trace: src/VX_lsu_mem_if.sv:5:15
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
										// Trace: src/VX_lsu_mem_if.sv:6:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_lsu_mem_if.sv:7:15
										localparam ADDR_WIDTH = 30;
										// Trace: src/VX_lsu_mem_if.sv:9:5
										localparam VX_gpu_pkg_UUID_WIDTH = 1;
										// removed localparam type tag_t
										// Trace: src/VX_lsu_mem_if.sv:13:5
										// removed localparam type req_data_t
										// Trace: src/VX_lsu_mem_if.sv:22:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_lsu_mem_if.sv:27:5
										wire req_valid;
										// Trace: src/VX_lsu_mem_if.sv:28:5
										wire [282:0] req_data;
										// Trace: src/VX_lsu_mem_if.sv:29:5
										wire req_ready;
										// Trace: src/VX_lsu_mem_if.sv:30:5
										wire rsp_valid;
										// Trace: src/VX_lsu_mem_if.sv:31:5
										wire [133:0] rsp_data;
										// Trace: src/VX_lsu_mem_if.sv:32:5
										wire rsp_ready;
										// Trace: src/VX_lsu_mem_if.sv:33:5
										// Trace: src/VX_lsu_mem_if.sv:41:5
									end
									// Trace: src/VX_mem_unit.sv:20:5
									genvar _gv_i_127;
									for (_gv_i_127 = 0; _gv_i_127 < 1; _gv_i_127 = _gv_i_127 + 1) begin : g_lmem_switches
										localparam i = _gv_i_127;
										// Trace: src/VX_mem_unit.sv:21:9
										// expanded module instance: lmem_switch
										localparam _bbase_5CF86_lsu_in_if = i + _mbase_lsu_mem_if;
										localparam _bbase_5CF86_global_out_if = i;
										localparam _bbase_5CF86_local_out_if = i;
										localparam _param_5CF86_GLOBAL_OUT_BUF = 1;
										localparam _param_5CF86_LOCAL_OUT_BUF = 1;
										localparam _param_5CF86_RSP_OUT_BUF = 1;
										localparam _param_5CF86_ARBITER = "P";
										if (1) begin : lmem_switch
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_lmem_switch.sv:2:15
											localparam GLOBAL_OUT_BUF = _param_5CF86_GLOBAL_OUT_BUF;
											// Trace: src/VX_lmem_switch.sv:3:15
											localparam LOCAL_OUT_BUF = _param_5CF86_LOCAL_OUT_BUF;
											// Trace: src/VX_lmem_switch.sv:4:15
											localparam RSP_OUT_BUF = _param_5CF86_RSP_OUT_BUF;
											// Trace: src/VX_lmem_switch.sv:5:15
											localparam ARBITER = _param_5CF86_ARBITER;
											// Trace: src/VX_lmem_switch.sv:7:5
											wire clk;
											// Trace: src/VX_lmem_switch.sv:8:5
											wire reset;
											// Trace: src/VX_lmem_switch.sv:9:5
											localparam _mbase_lsu_in_if = _bbase_5CF86_lsu_in_if;
											// Trace: src/VX_lmem_switch.sv:10:5
											localparam _mbase_global_out_if = _bbase_5CF86_global_out_if;
											// Trace: src/VX_lmem_switch.sv:11:5
											localparam _mbase_local_out_if = _bbase_5CF86_local_out_if;
											// Trace: src/VX_lmem_switch.sv:13:5
											localparam VX_gpu_pkg_XLENB = 4;
											localparam VX_gpu_pkg_LSU_WORD_SIZE = VX_gpu_pkg_XLENB;
											localparam VX_gpu_pkg_LSU_ADDR_WIDTH = 30;
											localparam VX_gpu_pkg_LSU_MEM_BATCHES = 1;
											localparam VX_gpu_pkg_LSU_TAG_ID_BITS = 1;
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											localparam VX_gpu_pkg_LSU_TAG_WIDTH = 2;
											localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
											localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
											localparam REQ_DATAW = 283;
											// Trace: src/VX_lmem_switch.sv:14:5
											localparam RSP_DATAW = 134;
											// Trace: src/VX_lmem_switch.sv:15:5
											wire [3:0] is_addr_local_mask;
											// Trace: src/VX_lmem_switch.sv:16:5
											wire req_global_ready;
											// Trace: src/VX_lmem_switch.sv:17:5
											wire req_local_ready;
											// Trace: src/VX_lmem_switch.sv:18:5
											genvar _gv_i_48;
											for (_gv_i_48 = 0; _gv_i_48 < 4; _gv_i_48 = _gv_i_48 + 1) begin : g_is_addr_local_mask
												localparam i = _gv_i_48;
												// Trace: src/VX_lmem_switch.sv:19:9
												assign is_addr_local_mask[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[2 + ((i * 3) + VX_gpu_pkg_MEM_REQ_FLAG_LOCAL)];
											end
											// Trace: src/VX_lmem_switch.sv:21:5
											wire is_addr_global = |(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[282-:4] & ~is_addr_local_mask);
											// Trace: src/VX_lmem_switch.sv:22:5
											wire is_addr_local = |(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[282-:4] & is_addr_local_mask);
											// Trace: src/VX_lmem_switch.sv:23:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_ready = (req_global_ready && is_addr_global) || (req_local_ready && is_addr_local);
											// Trace: src/VX_lmem_switch.sv:25:5
											VX_elastic_buffer #(
												.DATAW(REQ_DATAW),
												.SIZE(1),
												.OUT_REG(1)
											) req_global_buf(
												.clk(clk),
												.reset(reset),
												.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_valid && is_addr_global),
												.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[282-:4] & ~is_addr_local_mask, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[278], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[277-:120], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[157-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[29-:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[13-:12], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[1-:2]}),
												.ready_in(req_global_ready),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_dcache_if[_mbase_global_out_if].req_valid),
												.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_dcache_if[_mbase_global_out_if].req_data),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_dcache_if[_mbase_global_out_if].req_ready)
											);
											// Trace: src/VX_lmem_switch.sv:47:5
											VX_elastic_buffer #(
												.DATAW(REQ_DATAW),
												.SIZE(1),
												.OUT_REG(1)
											) req_local_buf(
												.clk(clk),
												.reset(reset),
												.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_valid && is_addr_local),
												.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[282-:4] & is_addr_local_mask, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[278], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[277-:120], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[157-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[29-:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[13-:12], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].req_data[1-:2]}),
												.ready_in(req_local_ready),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_local_out_if].req_valid),
												.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_local_out_if].req_data),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_local_out_if].req_ready)
											);
											// Trace: src/VX_lmem_switch.sv:69:5
											VX_stream_arb #(
												.NUM_INPUTS(2),
												.DATAW(RSP_DATAW),
												.ARBITER(ARBITER),
												.OUT_BUF(RSP_OUT_BUF)
											) rsp_arb(
												.clk(clk),
												.reset(reset),
												.valid_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_local_out_if].rsp_valid, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_dcache_if[_mbase_global_out_if].rsp_valid}),
												.ready_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_local_out_if].rsp_ready, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_dcache_if[_mbase_global_out_if].rsp_ready}),
												.data_in({Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[_mbase_local_out_if].rsp_data, Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_dcache_if[_mbase_global_out_if].rsp_data}),
												.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].rsp_data),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].rsp_valid),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.lsu_mem_if[_mbase_lsu_in_if].rsp_ready),
												.sel_out()
											);
										end
										assign lmem_switch.clk = clk;
										assign lmem_switch.reset = reset;
									end
									// Trace: src/VX_mem_unit.sv:34:5
									localparam VX_gpu_pkg_LMEM_TAG_WIDTH = 2;
									// expanded interface instance: lmem_arb_if
									localparam _param_CC10A_NUM_LANES = 4;
									localparam _param_CC10A_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
									localparam _param_CC10A_TAG_WIDTH = VX_gpu_pkg_LMEM_TAG_WIDTH;
									genvar _arr_CC10A;
									for (_arr_CC10A = 0; _arr_CC10A <= 0; _arr_CC10A = _arr_CC10A + 1) begin : lmem_arb_if
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_lsu_mem_if.sv:2:15
										localparam NUM_LANES = _param_CC10A_NUM_LANES;
										// Trace: src/VX_lsu_mem_if.sv:3:15
										localparam DATA_SIZE = _param_CC10A_DATA_SIZE;
										// Trace: src/VX_lsu_mem_if.sv:4:15
										localparam TAG_WIDTH = _param_CC10A_TAG_WIDTH;
										// Trace: src/VX_lsu_mem_if.sv:5:15
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
										// Trace: src/VX_lsu_mem_if.sv:6:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_lsu_mem_if.sv:7:15
										localparam ADDR_WIDTH = 30;
										// Trace: src/VX_lsu_mem_if.sv:9:5
										localparam VX_gpu_pkg_UUID_WIDTH = 1;
										// removed localparam type tag_t
										// Trace: src/VX_lsu_mem_if.sv:13:5
										// removed localparam type req_data_t
										// Trace: src/VX_lsu_mem_if.sv:22:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_lsu_mem_if.sv:27:5
										wire req_valid;
										// Trace: src/VX_lsu_mem_if.sv:28:5
										wire [282:0] req_data;
										// Trace: src/VX_lsu_mem_if.sv:29:5
										wire req_ready;
										// Trace: src/VX_lsu_mem_if.sv:30:5
										wire rsp_valid;
										// Trace: src/VX_lsu_mem_if.sv:31:5
										wire [133:0] rsp_data;
										// Trace: src/VX_lsu_mem_if.sv:32:5
										wire rsp_ready;
										// Trace: src/VX_lsu_mem_if.sv:33:5
										// Trace: src/VX_lsu_mem_if.sv:41:5
									end
									// Trace: src/VX_mem_unit.sv:39:5
									// expanded module instance: lmem_arb
									localparam _bbase_32A2E_bus_in_if = 0;
									localparam _bbase_32A2E_bus_out_if = 0;
									localparam _param_32A2E_NUM_INPUTS = 1;
									localparam _param_32A2E_NUM_OUTPUTS = 1;
									localparam _param_32A2E_NUM_LANES = 4;
									localparam _param_32A2E_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
									localparam _param_32A2E_TAG_WIDTH = VX_gpu_pkg_LSU_TAG_WIDTH;
									localparam _param_32A2E_TAG_SEL_IDX = 0;
									localparam _param_32A2E_ARBITER = "R";
									localparam _param_32A2E_REQ_OUT_BUF = 0;
									localparam _param_32A2E_RSP_OUT_BUF = 2;
									if (1) begin : lmem_arb
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_lsu_mem_arb.sv:2:15
										localparam NUM_INPUTS = _param_32A2E_NUM_INPUTS;
										// Trace: src/VX_lsu_mem_arb.sv:3:15
										localparam NUM_OUTPUTS = _param_32A2E_NUM_OUTPUTS;
										// Trace: src/VX_lsu_mem_arb.sv:4:15
										localparam NUM_LANES = _param_32A2E_NUM_LANES;
										// Trace: src/VX_lsu_mem_arb.sv:5:15
										localparam DATA_SIZE = _param_32A2E_DATA_SIZE;
										// Trace: src/VX_lsu_mem_arb.sv:6:15
										localparam TAG_WIDTH = _param_32A2E_TAG_WIDTH;
										// Trace: src/VX_lsu_mem_arb.sv:7:15
										localparam TAG_SEL_IDX = _param_32A2E_TAG_SEL_IDX;
										// Trace: src/VX_lsu_mem_arb.sv:8:15
										localparam REQ_OUT_BUF = _param_32A2E_REQ_OUT_BUF;
										// Trace: src/VX_lsu_mem_arb.sv:9:15
										localparam RSP_OUT_BUF = _param_32A2E_RSP_OUT_BUF;
										// Trace: src/VX_lsu_mem_arb.sv:10:15
										localparam ARBITER = _param_32A2E_ARBITER;
										// Trace: src/VX_lsu_mem_arb.sv:11:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_lsu_mem_arb.sv:12:15
										localparam ADDR_WIDTH = 30;
										// Trace: src/VX_lsu_mem_arb.sv:13:15
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
										// Trace: src/VX_lsu_mem_arb.sv:15:5
										wire clk;
										// Trace: src/VX_lsu_mem_arb.sv:16:5
										wire reset;
										// Trace: src/VX_lsu_mem_arb.sv:17:5
										localparam _mbase_bus_in_if = 0;
										// Trace: src/VX_lsu_mem_arb.sv:18:5
										localparam _mbase_bus_out_if = 0;
										// Trace: src/VX_lsu_mem_arb.sv:20:5
										localparam DATA_WIDTH = 32;
										// Trace: src/VX_lsu_mem_arb.sv:21:5
										localparam LOG_NUM_REQS = 0;
										// Trace: src/VX_lsu_mem_arb.sv:22:5
										localparam REQ_DATAW = 283;
										// Trace: src/VX_lsu_mem_arb.sv:23:5
										localparam RSP_DATAW = 134;
										// Trace: src/VX_lsu_mem_arb.sv:24:5
										wire [0:0] req_valid_out;
										// Trace: src/VX_lsu_mem_arb.sv:25:5
										wire [282:0] req_data_out;
										// Trace: src/VX_lsu_mem_arb.sv:26:5
										wire [0:0] req_ready_out;
										// Trace: src/VX_lsu_mem_arb.sv:27:5
										wire [0:0] req_sel_out;
										// Trace: src/VX_lsu_mem_arb.sv:28:5
										wire [0:0] req_valid_in;
										// Trace: src/VX_lsu_mem_arb.sv:29:5
										wire [282:0] req_data_in;
										// Trace: src/VX_lsu_mem_arb.sv:30:5
										wire [0:0] req_ready_in;
										// Trace: src/VX_lsu_mem_arb.sv:31:5
										genvar _gv_i_23;
										for (_gv_i_23 = 0; _gv_i_23 < NUM_INPUTS; _gv_i_23 = _gv_i_23 + 1) begin : g_req_data_in
											localparam i = _gv_i_23;
											// Trace: src/VX_lsu_mem_arb.sv:32:9
											assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[i + _mbase_bus_in_if].req_valid;
											// Trace: src/VX_lsu_mem_arb.sv:33:9
											assign req_data_in[i * 283+:283] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[i + _mbase_bus_in_if].req_data;
											// Trace: src/VX_lsu_mem_arb.sv:34:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[i + _mbase_bus_in_if].req_ready = req_ready_in[i];
										end
										// Trace: src/VX_lsu_mem_arb.sv:36:5
										VX_stream_arb #(
											.NUM_INPUTS(NUM_INPUTS),
											.NUM_OUTPUTS(NUM_OUTPUTS),
											.DATAW(REQ_DATAW),
											.ARBITER(ARBITER),
											.OUT_BUF(REQ_OUT_BUF)
										) req_arb(
											.clk(clk),
											.reset(reset),
											.valid_in(req_valid_in),
											.ready_in(req_ready_in),
											.data_in(req_data_in),
											.data_out(req_data_out),
											.sel_out(req_sel_out),
											.valid_out(req_valid_out),
											.ready_out(req_ready_out)
										);
										// Trace: src/VX_lsu_mem_arb.sv:53:5
										genvar _gv_i_24;
										for (_gv_i_24 = 0; _gv_i_24 < NUM_OUTPUTS; _gv_i_24 = _gv_i_24 + 1) begin : g_bus_out_if
											localparam i = _gv_i_24;
											// Trace: src/VX_lsu_mem_arb.sv:54:9
											wire [1:0] req_tag_out;
											// Trace: src/VX_lsu_mem_arb.sv:55:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[i + _mbase_bus_out_if].req_valid = req_valid_out[i];
											// Trace: src/VX_lsu_mem_arb.sv:56:9
											assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[i + _mbase_bus_out_if].req_data[282-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[i + _mbase_bus_out_if].req_data[278], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[i + _mbase_bus_out_if].req_data[277-:120], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[i + _mbase_bus_out_if].req_data[157-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[i + _mbase_bus_out_if].req_data[29-:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[i + _mbase_bus_out_if].req_data[13-:12], req_tag_out} = req_data_out[i * 283+:283];
											// Trace: src/VX_lsu_mem_arb.sv:65:9
											assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[i + _mbase_bus_out_if].req_ready;
											if (1) begin : g_req_tag_out
												// Trace: src/VX_lsu_mem_arb.sv:77:13
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[i + _mbase_bus_out_if].req_data[1-:2] = req_tag_out;
											end
										end
										// Trace: src/VX_lsu_mem_arb.sv:80:5
										wire [0:0] rsp_valid_out;
										// Trace: src/VX_lsu_mem_arb.sv:81:5
										wire [133:0] rsp_data_out;
										// Trace: src/VX_lsu_mem_arb.sv:82:5
										wire [0:0] rsp_ready_out;
										// Trace: src/VX_lsu_mem_arb.sv:83:5
										wire [0:0] rsp_valid_in;
										// Trace: src/VX_lsu_mem_arb.sv:84:5
										wire [133:0] rsp_data_in;
										// Trace: src/VX_lsu_mem_arb.sv:85:5
										wire [0:0] rsp_ready_in;
										// Trace: src/VX_lsu_mem_arb.sv:86:5
										if (1) begin : g_rsp_arb
											genvar _gv_i_26;
											for (_gv_i_26 = 0; _gv_i_26 < NUM_OUTPUTS; _gv_i_26 = _gv_i_26 + 1) begin : g_rsp_data_in
												localparam i = _gv_i_26;
												// Trace: src/VX_lsu_mem_arb.sv:125:13
												assign rsp_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[i + _mbase_bus_out_if].rsp_valid;
												// Trace: src/VX_lsu_mem_arb.sv:126:13
												assign rsp_data_in[i * 134+:134] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[i + _mbase_bus_out_if].rsp_data;
												// Trace: src/VX_lsu_mem_arb.sv:127:13
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[i + _mbase_bus_out_if].rsp_ready = rsp_ready_in[i];
											end
											// Trace: src/VX_lsu_mem_arb.sv:129:9
											VX_stream_arb #(
												.NUM_INPUTS(NUM_OUTPUTS),
												.NUM_OUTPUTS(NUM_INPUTS),
												.DATAW(RSP_DATAW),
												.ARBITER(ARBITER),
												.OUT_BUF(RSP_OUT_BUF)
											) req_arb(
												.clk(clk),
												.reset(reset),
												.valid_in(rsp_valid_in),
												.ready_in(rsp_ready_in),
												.data_in(rsp_data_in),
												.data_out(rsp_data_out),
												.valid_out(rsp_valid_out),
												.ready_out(rsp_ready_out),
												.sel_out()
											);
										end
										// Trace: src/VX_lsu_mem_arb.sv:147:5
										genvar _gv_i_27;
										for (_gv_i_27 = 0; _gv_i_27 < NUM_INPUTS; _gv_i_27 = _gv_i_27 + 1) begin : g_output
											localparam i = _gv_i_27;
											// Trace: src/VX_lsu_mem_arb.sv:148:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[i + _mbase_bus_in_if].rsp_valid = rsp_valid_out[i];
											// Trace: src/VX_lsu_mem_arb.sv:149:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[i + _mbase_bus_in_if].rsp_data = rsp_data_out[i * 134+:134];
											// Trace: src/VX_lsu_mem_arb.sv:150:9
											assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lsu_lmem_if[i + _mbase_bus_in_if].rsp_ready;
										end
									end
									assign lmem_arb.clk = clk;
									assign lmem_arb.reset = reset;
									// Trace: src/VX_mem_unit.sv:55:5
									// expanded interface instance: lmem_adapt_if
									localparam _param_8498F_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
									localparam _param_8498F_TAG_WIDTH = VX_gpu_pkg_LMEM_TAG_WIDTH;
									genvar _arr_8498F;
									for (_arr_8498F = 0; _arr_8498F <= 3; _arr_8498F = _arr_8498F + 1) begin : lmem_adapt_if
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_mem_bus_if.sv:2:15
										localparam DATA_SIZE = _param_8498F_DATA_SIZE;
										// Trace: src/VX_mem_bus_if.sv:3:15
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:4:15
										localparam TAG_WIDTH = _param_8498F_TAG_WIDTH;
										// Trace: src/VX_mem_bus_if.sv:5:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_mem_bus_if.sv:6:15
										localparam ADDR_WIDTH = 30;
										// Trace: src/VX_mem_bus_if.sv:8:5
										localparam VX_gpu_pkg_UUID_WIDTH = 1;
										// removed localparam type tag_t
										// Trace: src/VX_mem_bus_if.sv:12:5
										// removed localparam type req_data_t
										// Trace: src/VX_mem_bus_if.sv:20:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_mem_bus_if.sv:24:5
										wire req_valid;
										// Trace: src/VX_mem_bus_if.sv:25:5
										wire [71:0] req_data;
										// Trace: src/VX_mem_bus_if.sv:26:5
										wire req_ready;
										// Trace: src/VX_mem_bus_if.sv:27:5
										wire rsp_valid;
										// Trace: src/VX_mem_bus_if.sv:28:5
										wire [33:0] rsp_data;
										// Trace: src/VX_mem_bus_if.sv:29:5
										wire rsp_ready;
										// Trace: src/VX_mem_bus_if.sv:30:5
										// Trace: src/VX_mem_bus_if.sv:38:5
									end
									// Trace: src/VX_mem_unit.sv:59:5
									// expanded module instance: lmem_adapter
									localparam _bbase_ED918_lsu_mem_if = 0;
									localparam _bbase_ED918_mem_bus_if = 0;
									localparam _param_ED918_NUM_LANES = 4;
									localparam _param_ED918_DATA_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
									localparam _param_ED918_TAG_WIDTH = VX_gpu_pkg_LMEM_TAG_WIDTH;
									localparam _param_ED918_TAG_SEL_BITS = 1;
									localparam _param_ED918_ARBITER = "P";
									localparam _param_ED918_REQ_OUT_BUF = 3;
									localparam _param_ED918_RSP_OUT_BUF = 0;
									if (1) begin : lmem_adapter
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_lsu_adapter.sv:2:15
										localparam NUM_LANES = _param_ED918_NUM_LANES;
										// Trace: src/VX_lsu_adapter.sv:3:15
										localparam DATA_SIZE = _param_ED918_DATA_SIZE;
										// Trace: src/VX_lsu_adapter.sv:4:15
										localparam TAG_WIDTH = _param_ED918_TAG_WIDTH;
										// Trace: src/VX_lsu_adapter.sv:5:15
										localparam TAG_SEL_BITS = _param_ED918_TAG_SEL_BITS;
										// Trace: src/VX_lsu_adapter.sv:6:15
										localparam ARBITER = _param_ED918_ARBITER;
										// Trace: src/VX_lsu_adapter.sv:7:15
										localparam REQ_OUT_BUF = _param_ED918_REQ_OUT_BUF;
										// Trace: src/VX_lsu_adapter.sv:8:15
										localparam RSP_OUT_BUF = _param_ED918_RSP_OUT_BUF;
										// Trace: src/VX_lsu_adapter.sv:10:5
										wire clk;
										// Trace: src/VX_lsu_adapter.sv:11:5
										wire reset;
										// Trace: src/VX_lsu_adapter.sv:12:5
										localparam _mbase_lsu_mem_if = _bbase_ED918_lsu_mem_if;
										// Trace: src/VX_lsu_adapter.sv:13:5
										localparam _mbase_mem_bus_if = 0;
										// Trace: src/VX_lsu_adapter.sv:15:5
										localparam REQ_ADDR_WIDTH = 30;
										// Trace: src/VX_lsu_adapter.sv:16:5
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam REQ_DATA_WIDTH = 70;
										// Trace: src/VX_lsu_adapter.sv:17:5
										localparam RSP_DATA_WIDTH = 32;
										// Trace: src/VX_lsu_adapter.sv:18:5
										wire [279:0] req_data_in;
										// Trace: src/VX_lsu_adapter.sv:19:5
										wire [3:0] req_valid_out;
										// Trace: src/VX_lsu_adapter.sv:20:5
										wire [279:0] req_data_out;
										// Trace: src/VX_lsu_adapter.sv:21:5
										wire [7:0] req_tag_out;
										// Trace: src/VX_lsu_adapter.sv:22:5
										wire [3:0] req_ready_out;
										// Trace: src/VX_lsu_adapter.sv:23:5
										genvar _gv_i_177;
										for (_gv_i_177 = 0; _gv_i_177 < NUM_LANES; _gv_i_177 = _gv_i_177 + 1) begin : g_req_data_in
											localparam i = _gv_i_177;
											// Trace: src/VX_lsu_adapter.sv:24:9
											assign req_data_in[i * 70+:70] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].req_data[278], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].req_data[158 + (i * 30)+:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].req_data[30 + (i * 32)+:32], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].req_data[14 + (i * 4)+:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].req_data[2 + (i * 3)+:3]};
										end
										// Trace: src/VX_lsu_adapter.sv:32:5
										VX_stream_unpack #(
											.NUM_REQS(NUM_LANES),
											.DATA_WIDTH(REQ_DATA_WIDTH),
											.TAG_WIDTH(TAG_WIDTH),
											.OUT_BUF(REQ_OUT_BUF)
										) stream_unpack(
											.clk(clk),
											.reset(reset),
											.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].req_valid),
											.mask_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].req_data[282-:4]),
											.data_in(req_data_in),
											.tag_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].req_data[1-:2]),
											.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].req_ready),
											.valid_out(req_valid_out),
											.data_out(req_data_out),
											.tag_out(req_tag_out),
											.ready_out(req_ready_out)
										);
										// Trace: src/VX_lsu_adapter.sv:50:5
										genvar _gv_i_178;
										for (_gv_i_178 = 0; _gv_i_178 < NUM_LANES; _gv_i_178 = _gv_i_178 + 1) begin : g_mem_bus_req
											localparam i = _gv_i_178;
											// Trace: src/VX_lsu_adapter.sv:51:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_valid = req_valid_out[i];
											// Trace: src/VX_lsu_adapter.sv:52:9
											assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_data[71], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_data[70-:30], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_data[40-:32], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_data[8-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_data[4-:3]} = req_data_out[i * 70+:70];
											// Trace: src/VX_lsu_adapter.sv:59:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_data[1-:2] = req_tag_out[i * 2+:2];
											// Trace: src/VX_lsu_adapter.sv:60:9
											assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_ready;
										end
										// Trace: src/VX_lsu_adapter.sv:62:5
										wire [3:0] rsp_valid_out;
										// Trace: src/VX_lsu_adapter.sv:63:5
										wire [127:0] rsp_data_out;
										// Trace: src/VX_lsu_adapter.sv:64:5
										wire [7:0] rsp_tag_out;
										// Trace: src/VX_lsu_adapter.sv:65:5
										wire [3:0] rsp_ready_out;
										// Trace: src/VX_lsu_adapter.sv:66:5
										genvar _gv_i_179;
										for (_gv_i_179 = 0; _gv_i_179 < NUM_LANES; _gv_i_179 = _gv_i_179 + 1) begin : g_mem_bus_rsp
											localparam i = _gv_i_179;
											// Trace: src/VX_lsu_adapter.sv:67:9
											assign rsp_valid_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].rsp_valid;
											// Trace: src/VX_lsu_adapter.sv:68:9
											assign rsp_data_out[i * 32+:32] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].rsp_data[33-:32];
											// Trace: src/VX_lsu_adapter.sv:69:9
											assign rsp_tag_out[i * 2+:2] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].rsp_data[1-:2];
											// Trace: src/VX_lsu_adapter.sv:70:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].rsp_ready = rsp_ready_out[i];
										end
										// Trace: src/VX_lsu_adapter.sv:72:5
										VX_stream_pack #(
											.NUM_REQS(NUM_LANES),
											.DATA_WIDTH(RSP_DATA_WIDTH),
											.TAG_WIDTH(TAG_WIDTH),
											.TAG_SEL_BITS(TAG_SEL_BITS),
											.ARBITER(ARBITER),
											.OUT_BUF(RSP_OUT_BUF)
										) stream_pack(
											.clk(clk),
											.reset(reset),
											.valid_in(rsp_valid_out),
											.data_in(rsp_data_out),
											.tag_in(rsp_tag_out),
											.ready_in(rsp_ready_out),
											.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].rsp_valid),
											.mask_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].rsp_data[133-:4]),
											.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].rsp_data[129-:128]),
											.tag_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].rsp_data[1-:2]),
											.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_arb_if[_mbase_lsu_mem_if].rsp_ready)
										);
									end
									assign lmem_adapter.clk = clk;
									assign lmem_adapter.reset = reset;
									// Trace: src/VX_mem_unit.sv:73:5
									// expanded module instance: local_mem
									localparam _bbase_9EDEE_mem_bus_if = 0;
									localparam _param_9EDEE_INSTANCE_ID = "";
									localparam _param_9EDEE_SIZE = 16384;
									localparam _param_9EDEE_NUM_REQS = 4;
									localparam _param_9EDEE_NUM_BANKS = 4;
									localparam _param_9EDEE_WORD_SIZE = VX_gpu_pkg_LSU_WORD_SIZE;
									localparam _param_9EDEE_ADDR_WIDTH = LMEM_ADDR_WIDTH;
									localparam _param_9EDEE_TAG_WIDTH = VX_gpu_pkg_LMEM_TAG_WIDTH;
									localparam _param_9EDEE_OUT_BUF = 3;
									if (1) begin : local_mem
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_local_mem.sv:2:15
										localparam INSTANCE_ID = _param_9EDEE_INSTANCE_ID;
										// Trace: src/VX_local_mem.sv:3:15
										localparam SIZE = _param_9EDEE_SIZE;
										// Trace: src/VX_local_mem.sv:4:15
										localparam NUM_REQS = _param_9EDEE_NUM_REQS;
										// Trace: src/VX_local_mem.sv:5:15
										localparam NUM_BANKS = _param_9EDEE_NUM_BANKS;
										// Trace: src/VX_local_mem.sv:6:15
										localparam ADDR_WIDTH = _param_9EDEE_ADDR_WIDTH;
										// Trace: src/VX_local_mem.sv:7:15
										localparam WORD_SIZE = _param_9EDEE_WORD_SIZE;
										// Trace: src/VX_local_mem.sv:8:15
										localparam TAG_WIDTH = _param_9EDEE_TAG_WIDTH;
										// Trace: src/VX_local_mem.sv:9:15
										localparam OUT_BUF = _param_9EDEE_OUT_BUF;
										// Trace: src/VX_local_mem.sv:11:5
										wire clk;
										// Trace: src/VX_local_mem.sv:12:5
										wire reset;
										// Trace: src/VX_local_mem.sv:13:5
										localparam _mbase_mem_bus_if = 0;
										// Trace: src/VX_local_mem.sv:15:5
										localparam REQ_SEL_BITS = 2;
										// Trace: src/VX_local_mem.sv:16:5
										localparam REQ_SEL_WIDTH = REQ_SEL_BITS;
										// Trace: src/VX_local_mem.sv:17:5
										localparam WORD_WIDTH = 32;
										// Trace: src/VX_local_mem.sv:18:5
										localparam NUM_WORDS = 4096;
										// Trace: src/VX_local_mem.sv:19:5
										localparam WORDS_PER_BANK = 1024;
										// Trace: src/VX_local_mem.sv:20:5
										localparam BANK_ADDR_WIDTH = 10;
										// Trace: src/VX_local_mem.sv:21:5
										localparam BANK_SEL_BITS = 2;
										// Trace: src/VX_local_mem.sv:22:5
										localparam BANK_SEL_WIDTH = BANK_SEL_BITS;
										// Trace: src/VX_local_mem.sv:23:5
										localparam REQ_DATAW = 49;
										// Trace: src/VX_local_mem.sv:24:5
										localparam RSP_DATAW = 34;
										// Trace: src/VX_local_mem.sv:25:5
										wire [7:0] req_bank_idx;
										// Trace: src/VX_local_mem.sv:26:5
										if (1) begin : g_req_bank_idx
											genvar _gv_i_196;
											for (_gv_i_196 = 0; _gv_i_196 < NUM_REQS; _gv_i_196 = _gv_i_196 + 1) begin : g_req_bank_idxs
												localparam i = _gv_i_196;
												// Trace: src/VX_local_mem.sv:28:13
												assign req_bank_idx[i * 2+:2] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_data[41+:BANK_SEL_BITS];
											end
										end
										// Trace: src/VX_local_mem.sv:33:5
										wire [39:0] req_bank_addr;
										// Trace: src/VX_local_mem.sv:34:5
										genvar _gv_i_197;
										for (_gv_i_197 = 0; _gv_i_197 < NUM_REQS; _gv_i_197 = _gv_i_197 + 1) begin : g_req_bank_addr
											localparam i = _gv_i_197;
											// Trace: src/VX_local_mem.sv:35:9
											assign req_bank_addr[i * 10+:10] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_data[43+:BANK_ADDR_WIDTH];
										end
										// Trace: src/VX_local_mem.sv:37:5
										wire [3:0] per_bank_req_valid;
										// Trace: src/VX_local_mem.sv:38:5
										wire [3:0] per_bank_req_rw;
										// Trace: src/VX_local_mem.sv:39:5
										wire [39:0] per_bank_req_addr;
										// Trace: src/VX_local_mem.sv:40:5
										wire [15:0] per_bank_req_byteen;
										// Trace: src/VX_local_mem.sv:41:5
										wire [127:0] per_bank_req_data;
										// Trace: src/VX_local_mem.sv:42:5
										wire [7:0] per_bank_req_tag;
										// Trace: src/VX_local_mem.sv:43:5
										wire [7:0] per_bank_req_idx;
										// Trace: src/VX_local_mem.sv:44:5
										wire [3:0] per_bank_req_ready;
										// Trace: src/VX_local_mem.sv:45:5
										wire [195:0] per_bank_req_data_aos;
										// Trace: src/VX_local_mem.sv:46:5
										wire [3:0] req_valid_in;
										// Trace: src/VX_local_mem.sv:47:5
										wire [195:0] req_data_in;
										// Trace: src/VX_local_mem.sv:48:5
										wire [3:0] req_ready_in;
										// Trace: src/VX_local_mem.sv:49:5
										genvar _gv_i_198;
										for (_gv_i_198 = 0; _gv_i_198 < NUM_REQS; _gv_i_198 = _gv_i_198 + 1) begin : g_req_data_in
											localparam i = _gv_i_198;
											// Trace: src/VX_local_mem.sv:50:9
											assign req_valid_in[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_valid;
											// Trace: src/VX_local_mem.sv:51:9
											assign req_data_in[i * 49+:49] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_data[71], req_bank_addr[i * 10+:10], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_data[40-:32], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_data[8-:4], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_data[1-:2]};
											// Trace: src/VX_local_mem.sv:58:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].req_ready = req_ready_in[i];
										end
										// Trace: src/VX_local_mem.sv:60:5
										localparam VX_gpu_pkg_PERF_CTR_BITS = 44;
										VX_stream_xbar #(
											.NUM_INPUTS(NUM_REQS),
											.NUM_OUTPUTS(NUM_BANKS),
											.DATAW(REQ_DATAW),
											.PERF_CTR_BITS(VX_gpu_pkg_PERF_CTR_BITS),
											.ARBITER("P"),
											.OUT_BUF(3)
										) req_xbar(
											.clk(clk),
											.reset(reset),
											.collisions(),
											.valid_in(req_valid_in),
											.data_in(req_data_in),
											.sel_in(req_bank_idx),
											.ready_in(req_ready_in),
											.valid_out(per_bank_req_valid),
											.data_out(per_bank_req_data_aos),
											.sel_out(per_bank_req_idx),
											.ready_out(per_bank_req_ready)
										);
										// Trace: src/VX_local_mem.sv:80:5
										genvar _gv_i_199;
										for (_gv_i_199 = 0; _gv_i_199 < NUM_BANKS; _gv_i_199 = _gv_i_199 + 1) begin : g_per_bank_req_data_soa
											localparam i = _gv_i_199;
											// Trace: src/VX_local_mem.sv:81:9
											assign {per_bank_req_rw[i], per_bank_req_addr[i * 10+:10], per_bank_req_data[i * 32+:32], per_bank_req_byteen[i * 4+:4], per_bank_req_tag[i * 2+:2]} = per_bank_req_data_aos[i * 49+:49];
										end
										// Trace: src/VX_local_mem.sv:89:5
										wire [3:0] per_bank_rsp_valid;
										// Trace: src/VX_local_mem.sv:90:5
										wire [127:0] per_bank_rsp_data;
										// Trace: src/VX_local_mem.sv:91:5
										wire [7:0] per_bank_rsp_idx;
										// Trace: src/VX_local_mem.sv:92:5
										wire [7:0] per_bank_rsp_tag;
										// Trace: src/VX_local_mem.sv:93:5
										wire [3:0] per_bank_rsp_ready;
										// Trace: src/VX_local_mem.sv:94:5
										genvar _gv_i_200;
										for (_gv_i_200 = 0; _gv_i_200 < NUM_BANKS; _gv_i_200 = _gv_i_200 + 1) begin : g_data_store
											localparam i = _gv_i_200;
											// Trace: src/VX_local_mem.sv:95:9
											wire bank_rsp_valid;
											wire bank_rsp_ready;
											// Trace: src/VX_local_mem.sv:96:9
											VX_sp_ram #(
												.DATAW(WORD_WIDTH),
												.SIZE(WORDS_PER_BANK),
												.WRENW(WORD_SIZE),
												.OUT_REG(1),
												.RDW_MODE("R")
											) lmem_store(
												.clk(clk),
												.reset(reset),
												.read((per_bank_req_valid[i] && per_bank_req_ready[i]) && ~per_bank_req_rw[i]),
												.write((per_bank_req_valid[i] && per_bank_req_ready[i]) && per_bank_req_rw[i]),
												.wren(per_bank_req_byteen[i * 4+:4]),
												.addr(per_bank_req_addr[i * 10+:10]),
												.wdata(per_bank_req_data[i * 32+:32]),
												.rdata(per_bank_rsp_data[i * 32+:32])
											);
											// Trace: src/VX_local_mem.sv:112:9
											reg [9:0] last_wr_addr;
											// Trace: src/VX_local_mem.sv:113:9
											reg last_wr_valid;
											// Trace: src/VX_local_mem.sv:114:9
											always @(posedge clk) begin
												// Trace: src/VX_local_mem.sv:115:13
												if (reset)
													// Trace: src/VX_local_mem.sv:116:17
													last_wr_valid <= 0;
												else
													// Trace: src/VX_local_mem.sv:118:17
													last_wr_valid <= (per_bank_req_valid[i] && per_bank_req_ready[i]) && per_bank_req_rw[i];
												// Trace: src/VX_local_mem.sv:120:13
												last_wr_addr <= per_bank_req_addr[i * 10+:10];
											end
											// Trace: src/VX_local_mem.sv:122:9
											wire is_rdw_hazard = (last_wr_valid && ~per_bank_req_rw[i]) && (per_bank_req_addr[i * 10+:10] == last_wr_addr);
											// Trace: src/VX_local_mem.sv:123:9
											assign bank_rsp_valid = (per_bank_req_valid[i] && ~per_bank_req_rw[i]) && ~is_rdw_hazard;
											// Trace: src/VX_local_mem.sv:124:9
											assign per_bank_req_ready[i] = (bank_rsp_ready || per_bank_req_rw[i]) && ~is_rdw_hazard;
											// Trace: src/VX_local_mem.sv:125:9
											VX_pipe_buffer #(.DATAW(4)) bram_buf(
												.clk(clk),
												.reset(reset),
												.valid_in(bank_rsp_valid),
												.ready_in(bank_rsp_ready),
												.data_in({per_bank_req_idx[i * 2+:2], per_bank_req_tag[i * 2+:2]}),
												.data_out({per_bank_rsp_idx[i * 2+:2], per_bank_rsp_tag[i * 2+:2]}),
												.valid_out(per_bank_rsp_valid[i]),
												.ready_out(per_bank_rsp_ready[i])
											);
										end
										// Trace: src/VX_local_mem.sv:138:5
										wire [135:0] per_bank_rsp_data_aos;
										// Trace: src/VX_local_mem.sv:139:5
										genvar _gv_i_201;
										for (_gv_i_201 = 0; _gv_i_201 < NUM_BANKS; _gv_i_201 = _gv_i_201 + 1) begin : g_per_bank_rsp_data_aos
											localparam i = _gv_i_201;
											// Trace: src/VX_local_mem.sv:140:9
											assign per_bank_rsp_data_aos[i * 34+:34] = {per_bank_rsp_data[i * 32+:32], per_bank_rsp_tag[i * 2+:2]};
										end
										// Trace: src/VX_local_mem.sv:142:5
										wire [3:0] rsp_valid_out;
										// Trace: src/VX_local_mem.sv:143:5
										wire [135:0] rsp_data_out;
										// Trace: src/VX_local_mem.sv:144:5
										wire [3:0] rsp_ready_out;
										// Trace: src/VX_local_mem.sv:145:5
										VX_stream_xbar #(
											.NUM_INPUTS(NUM_BANKS),
											.NUM_OUTPUTS(NUM_REQS),
											.DATAW(RSP_DATAW),
											.ARBITER("P"),
											.OUT_BUF(OUT_BUF)
										) rsp_xbar(
											.clk(clk),
											.reset(reset),
											.collisions(),
											.sel_in(per_bank_rsp_idx),
											.valid_in(per_bank_rsp_valid),
											.data_in(per_bank_rsp_data_aos),
											.ready_in(per_bank_rsp_ready),
											.valid_out(rsp_valid_out),
											.data_out(rsp_data_out),
											.ready_out(rsp_ready_out),
											.sel_out()
										);
										// Trace: src/VX_local_mem.sv:164:5
										genvar _gv_i_202;
										for (_gv_i_202 = 0; _gv_i_202 < NUM_REQS; _gv_i_202 = _gv_i_202 + 1) begin : g_mem_bus_if
											localparam i = _gv_i_202;
											// Trace: src/VX_local_mem.sv:165:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].rsp_valid = rsp_valid_out[i];
											// Trace: src/VX_local_mem.sv:166:9
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].rsp_data = rsp_data_out[i * 34+:34];
											// Trace: src/VX_local_mem.sv:167:9
											assign rsp_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.lmem_adapt_if[i + _mbase_mem_bus_if].rsp_ready;
										end
									end
									assign local_mem.clk = clk;
									assign local_mem.reset = reset;
									// Trace: src/VX_mem_unit.sv:87:5
									localparam VX_gpu_pkg_DCACHE_MERGED_REQS = 1;
									localparam VX_gpu_pkg_DCACHE_MEM_BATCHES = 1;
									localparam VX_gpu_pkg_DCACHE_TAG_ID_BITS = 2;
									localparam VX_gpu_pkg_DCACHE_TAG_WIDTH = 3;
									// expanded interface instance: dcache_coalesced_if
									localparam _param_419A9_NUM_LANES = VX_gpu_pkg_DCACHE_CHANNELS;
									localparam _param_419A9_DATA_SIZE = VX_gpu_pkg_DCACHE_WORD_SIZE;
									localparam _param_419A9_TAG_WIDTH = VX_gpu_pkg_DCACHE_TAG_WIDTH;
									genvar _arr_419A9;
									for (_arr_419A9 = 0; _arr_419A9 <= 0; _arr_419A9 = _arr_419A9 + 1) begin : dcache_coalesced_if
										// removed import VX_gpu_pkg::*;
										// Trace: src/VX_lsu_mem_if.sv:2:15
										localparam NUM_LANES = _param_419A9_NUM_LANES;
										// Trace: src/VX_lsu_mem_if.sv:3:15
										localparam DATA_SIZE = _param_419A9_DATA_SIZE;
										// Trace: src/VX_lsu_mem_if.sv:4:15
										localparam TAG_WIDTH = _param_419A9_TAG_WIDTH;
										// Trace: src/VX_lsu_mem_if.sv:5:15
										localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
										localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
										localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
										// Trace: src/VX_lsu_mem_if.sv:6:15
										localparam MEM_ADDR_WIDTH = 32;
										// Trace: src/VX_lsu_mem_if.sv:7:15
										localparam ADDR_WIDTH = 28;
										// Trace: src/VX_lsu_mem_if.sv:9:5
										localparam VX_gpu_pkg_UUID_WIDTH = 1;
										// removed localparam type tag_t
										// Trace: src/VX_lsu_mem_if.sv:13:5
										// removed localparam type req_data_t
										// Trace: src/VX_lsu_mem_if.sv:22:5
										// removed localparam type rsp_data_t
										// Trace: src/VX_lsu_mem_if.sv:27:5
										wire req_valid;
										// Trace: src/VX_lsu_mem_if.sv:28:5
										wire [179:0] req_data;
										// Trace: src/VX_lsu_mem_if.sv:29:5
										wire req_ready;
										// Trace: src/VX_lsu_mem_if.sv:30:5
										wire rsp_valid;
										// Trace: src/VX_lsu_mem_if.sv:31:5
										wire [131:0] rsp_data;
										// Trace: src/VX_lsu_mem_if.sv:32:5
										wire rsp_ready;
										// Trace: src/VX_lsu_mem_if.sv:33:5
										// Trace: src/VX_lsu_mem_if.sv:41:5
									end
									// Trace: src/VX_mem_unit.sv:92:5
									localparam VX_gpu_pkg_LSU_ADDR_WIDTH = 30;
									localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
									localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
									localparam VX_gpu_pkg_PERF_CTR_BITS = 44;
									if (1) begin : g_enabled
										genvar _gv_i_128;
										for (_gv_i_128 = 0; _gv_i_128 < 1; _gv_i_128 = _gv_i_128 + 1) begin : g_coalescers
											localparam i = _gv_i_128;
											// Trace: src/VX_mem_unit.sv:94:13
											VX_mem_coalescer #(
												.INSTANCE_ID(""),
												.NUM_REQS(4),
												.DATA_IN_SIZE(VX_gpu_pkg_LSU_WORD_SIZE),
												.DATA_OUT_SIZE(VX_gpu_pkg_DCACHE_WORD_SIZE),
												.ADDR_WIDTH(VX_gpu_pkg_LSU_ADDR_WIDTH),
												.FLAGS_WIDTH(VX_gpu_pkg_MEM_FLAGS_WIDTH),
												.TAG_WIDTH(VX_gpu_pkg_LSU_TAG_WIDTH),
												.UUID_WIDTH(VX_gpu_pkg_UUID_WIDTH),
												.QUEUE_SIZE(4),
												.PERF_CTR_BITS(VX_gpu_pkg_PERF_CTR_BITS)
											) mem_coalescer(
												.clk(clk),
												.reset(reset),
												.misses(),
												.in_req_valid(lsu_dcache_if[i].req_valid),
												.in_req_mask(lsu_dcache_if[i].req_data[282-:4]),
												.in_req_rw(lsu_dcache_if[i].req_data[278]),
												.in_req_byteen(lsu_dcache_if[i].req_data[29-:16]),
												.in_req_addr(lsu_dcache_if[i].req_data[277-:120]),
												.in_req_flags(lsu_dcache_if[i].req_data[13-:12]),
												.in_req_data(lsu_dcache_if[i].req_data[157-:128]),
												.in_req_tag(lsu_dcache_if[i].req_data[1-:2]),
												.in_req_ready(lsu_dcache_if[i].req_ready),
												.in_rsp_valid(lsu_dcache_if[i].rsp_valid),
												.in_rsp_mask(lsu_dcache_if[i].rsp_data[133-:4]),
												.in_rsp_data(lsu_dcache_if[i].rsp_data[129-:128]),
												.in_rsp_tag(lsu_dcache_if[i].rsp_data[1-:2]),
												.in_rsp_ready(lsu_dcache_if[i].rsp_ready),
												.out_req_valid(dcache_coalesced_if[i].req_valid),
												.out_req_mask(dcache_coalesced_if[i].req_data[179-:1]),
												.out_req_rw(dcache_coalesced_if[i].req_data[178]),
												.out_req_byteen(dcache_coalesced_if[i].req_data[21-:16]),
												.out_req_addr(dcache_coalesced_if[i].req_data[177-:28]),
												.out_req_flags(dcache_coalesced_if[i].req_data[5-:3]),
												.out_req_data(dcache_coalesced_if[i].req_data[149-:128]),
												.out_req_tag(dcache_coalesced_if[i].req_data[2-:3]),
												.out_req_ready(dcache_coalesced_if[i].req_ready),
												.out_rsp_valid(dcache_coalesced_if[i].rsp_valid),
												.out_rsp_mask(dcache_coalesced_if[i].rsp_data[131-:1]),
												.out_rsp_data(dcache_coalesced_if[i].rsp_data[130-:128]),
												.out_rsp_tag(dcache_coalesced_if[i].rsp_data[2-:3]),
												.out_rsp_ready(dcache_coalesced_if[i].rsp_ready)
											);
										end
									end
									// Trace: src/VX_mem_unit.sv:149:5
									genvar _gv_i_130;
									for (_gv_i_130 = 0; _gv_i_130 < 1; _gv_i_130 = _gv_i_130 + 1) begin : g_dcache_adapters
										localparam i = _gv_i_130;
										// Trace: src/VX_mem_unit.sv:150:9
										// expanded interface instance: dcache_bus_tmp_if
										localparam _param_CE5A6_DATA_SIZE = VX_gpu_pkg_DCACHE_WORD_SIZE;
										localparam _param_CE5A6_TAG_WIDTH = VX_gpu_pkg_DCACHE_TAG_WIDTH;
										genvar _arr_CE5A6;
										for (_arr_CE5A6 = 0; _arr_CE5A6 <= 0; _arr_CE5A6 = _arr_CE5A6 + 1) begin : dcache_bus_tmp_if
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_mem_bus_if.sv:2:15
											localparam DATA_SIZE = _param_CE5A6_DATA_SIZE;
											// Trace: src/VX_mem_bus_if.sv:3:15
											localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
											localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
											localparam FLAGS_WIDTH = VX_gpu_pkg_MEM_FLAGS_WIDTH;
											// Trace: src/VX_mem_bus_if.sv:4:15
											localparam TAG_WIDTH = _param_CE5A6_TAG_WIDTH;
											// Trace: src/VX_mem_bus_if.sv:5:15
											localparam MEM_ADDR_WIDTH = 32;
											// Trace: src/VX_mem_bus_if.sv:6:15
											localparam ADDR_WIDTH = 28;
											// Trace: src/VX_mem_bus_if.sv:8:5
											localparam VX_gpu_pkg_UUID_WIDTH = 1;
											// removed localparam type tag_t
											// Trace: src/VX_mem_bus_if.sv:12:5
											// removed localparam type req_data_t
											// Trace: src/VX_mem_bus_if.sv:20:5
											// removed localparam type rsp_data_t
											// Trace: src/VX_mem_bus_if.sv:24:5
											wire req_valid;
											// Trace: src/VX_mem_bus_if.sv:25:5
											wire [178:0] req_data;
											// Trace: src/VX_mem_bus_if.sv:26:5
											wire req_ready;
											// Trace: src/VX_mem_bus_if.sv:27:5
											wire rsp_valid;
											// Trace: src/VX_mem_bus_if.sv:28:5
											wire [130:0] rsp_data;
											// Trace: src/VX_mem_bus_if.sv:29:5
											wire rsp_ready;
											// Trace: src/VX_mem_bus_if.sv:30:5
											// Trace: src/VX_mem_bus_if.sv:38:5
										end
										// Trace: src/VX_mem_unit.sv:154:9
										// expanded module instance: dcache_adapter
										localparam _bbase_6EE01_lsu_mem_if = i;
										localparam _bbase_6EE01_mem_bus_if = 0;
										localparam _param_6EE01_NUM_LANES = VX_gpu_pkg_DCACHE_CHANNELS;
										localparam _param_6EE01_DATA_SIZE = VX_gpu_pkg_DCACHE_WORD_SIZE;
										localparam _param_6EE01_TAG_WIDTH = VX_gpu_pkg_DCACHE_TAG_WIDTH;
										localparam _param_6EE01_TAG_SEL_BITS = 2;
										localparam _param_6EE01_ARBITER = "P";
										localparam _param_6EE01_REQ_OUT_BUF = 0;
										localparam _param_6EE01_RSP_OUT_BUF = 0;
										if (1) begin : dcache_adapter
											// removed import VX_gpu_pkg::*;
											// Trace: src/VX_lsu_adapter.sv:2:15
											localparam NUM_LANES = _param_6EE01_NUM_LANES;
											// Trace: src/VX_lsu_adapter.sv:3:15
											localparam DATA_SIZE = _param_6EE01_DATA_SIZE;
											// Trace: src/VX_lsu_adapter.sv:4:15
											localparam TAG_WIDTH = _param_6EE01_TAG_WIDTH;
											// Trace: src/VX_lsu_adapter.sv:5:15
											localparam TAG_SEL_BITS = _param_6EE01_TAG_SEL_BITS;
											// Trace: src/VX_lsu_adapter.sv:6:15
											localparam ARBITER = _param_6EE01_ARBITER;
											// Trace: src/VX_lsu_adapter.sv:7:15
											localparam REQ_OUT_BUF = _param_6EE01_REQ_OUT_BUF;
											// Trace: src/VX_lsu_adapter.sv:8:15
											localparam RSP_OUT_BUF = _param_6EE01_RSP_OUT_BUF;
											// Trace: src/VX_lsu_adapter.sv:10:5
											wire clk;
											// Trace: src/VX_lsu_adapter.sv:11:5
											wire reset;
											// Trace: src/VX_lsu_adapter.sv:12:5
											localparam _mbase_lsu_mem_if = _bbase_6EE01_lsu_mem_if;
											// Trace: src/VX_lsu_adapter.sv:13:5
											localparam _mbase_mem_bus_if = 0;
											// Trace: src/VX_lsu_adapter.sv:15:5
											localparam REQ_ADDR_WIDTH = 28;
											// Trace: src/VX_lsu_adapter.sv:16:5
											localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
											localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
											localparam REQ_DATA_WIDTH = 176;
											// Trace: src/VX_lsu_adapter.sv:17:5
											localparam RSP_DATA_WIDTH = 128;
											// Trace: src/VX_lsu_adapter.sv:18:5
											wire [175:0] req_data_in;
											// Trace: src/VX_lsu_adapter.sv:19:5
											wire [0:0] req_valid_out;
											// Trace: src/VX_lsu_adapter.sv:20:5
											wire [175:0] req_data_out;
											// Trace: src/VX_lsu_adapter.sv:21:5
											wire [2:0] req_tag_out;
											// Trace: src/VX_lsu_adapter.sv:22:5
											wire [0:0] req_ready_out;
											// Trace: src/VX_lsu_adapter.sv:23:5
											genvar _gv_i_177;
											for (_gv_i_177 = 0; _gv_i_177 < NUM_LANES; _gv_i_177 = _gv_i_177 + 1) begin : g_req_data_in
												localparam i = _gv_i_177;
												// Trace: src/VX_lsu_adapter.sv:24:9
												assign req_data_in[i * 176+:176] = {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[178], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[150 + (i * 28)+:28], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[22 + (i * 128)+:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[6 + (i * 16)+:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[3 + (i * 3)+:3]};
											end
											// Trace: src/VX_lsu_adapter.sv:32:5
											VX_stream_unpack #(
												.NUM_REQS(NUM_LANES),
												.DATA_WIDTH(REQ_DATA_WIDTH),
												.TAG_WIDTH(TAG_WIDTH),
												.OUT_BUF(REQ_OUT_BUF)
											) stream_unpack(
												.clk(clk),
												.reset(reset),
												.valid_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_valid),
												.mask_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[179-:1]),
												.data_in(req_data_in),
												.tag_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_data[2-:3]),
												.ready_in(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].req_ready),
												.valid_out(req_valid_out),
												.data_out(req_data_out),
												.tag_out(req_tag_out),
												.ready_out(req_ready_out)
											);
											// Trace: src/VX_lsu_adapter.sv:50:5
											genvar _gv_i_178;
											for (_gv_i_178 = 0; _gv_i_178 < NUM_LANES; _gv_i_178 = _gv_i_178 + 1) begin : g_mem_bus_req
												localparam i = _gv_i_178;
												// Trace: src/VX_lsu_adapter.sv:51:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_130].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_valid = req_valid_out[i];
												// Trace: src/VX_lsu_adapter.sv:52:9
												assign {Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_130].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_data[178], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_130].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_data[177-:28], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_130].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_data[149-:128], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_130].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_data[21-:16], Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_130].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_data[5-:3]} = req_data_out[i * 176+:176];
												// Trace: src/VX_lsu_adapter.sv:59:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_130].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_data[2-:3] = req_tag_out[i * 3+:3];
												// Trace: src/VX_lsu_adapter.sv:60:9
												assign req_ready_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_130].dcache_bus_tmp_if[i + _mbase_mem_bus_if].req_ready;
											end
											// Trace: src/VX_lsu_adapter.sv:62:5
											wire [0:0] rsp_valid_out;
											// Trace: src/VX_lsu_adapter.sv:63:5
											wire [127:0] rsp_data_out;
											// Trace: src/VX_lsu_adapter.sv:64:5
											wire [2:0] rsp_tag_out;
											// Trace: src/VX_lsu_adapter.sv:65:5
											wire [0:0] rsp_ready_out;
											// Trace: src/VX_lsu_adapter.sv:66:5
											genvar _gv_i_179;
											for (_gv_i_179 = 0; _gv_i_179 < NUM_LANES; _gv_i_179 = _gv_i_179 + 1) begin : g_mem_bus_rsp
												localparam i = _gv_i_179;
												// Trace: src/VX_lsu_adapter.sv:67:9
												assign rsp_valid_out[i] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_130].dcache_bus_tmp_if[i + _mbase_mem_bus_if].rsp_valid;
												// Trace: src/VX_lsu_adapter.sv:68:9
												assign rsp_data_out[i * 128+:128] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_130].dcache_bus_tmp_if[i + _mbase_mem_bus_if].rsp_data[130-:128];
												// Trace: src/VX_lsu_adapter.sv:69:9
												assign rsp_tag_out[i * 3+:3] = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_130].dcache_bus_tmp_if[i + _mbase_mem_bus_if].rsp_data[2-:3];
												// Trace: src/VX_lsu_adapter.sv:70:9
												assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.g_dcache_adapters[_gv_i_130].dcache_bus_tmp_if[i + _mbase_mem_bus_if].rsp_ready = rsp_ready_out[i];
											end
											// Trace: src/VX_lsu_adapter.sv:72:5
											VX_stream_pack #(
												.NUM_REQS(NUM_LANES),
												.DATA_WIDTH(RSP_DATA_WIDTH),
												.TAG_WIDTH(TAG_WIDTH),
												.TAG_SEL_BITS(TAG_SEL_BITS),
												.ARBITER(ARBITER),
												.OUT_BUF(RSP_OUT_BUF)
											) stream_pack(
												.clk(clk),
												.reset(reset),
												.valid_in(rsp_valid_out),
												.data_in(rsp_data_out),
												.tag_in(rsp_tag_out),
												.ready_in(rsp_ready_out),
												.valid_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].rsp_valid),
												.mask_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].rsp_data[131-:1]),
												.data_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].rsp_data[130-:128]),
												.tag_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].rsp_data[2-:3]),
												.ready_out(Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.g_cores[_gv_core_id_1].core.mem_unit.dcache_coalesced_if[_mbase_lsu_mem_if].rsp_ready)
											);
										end
										assign dcache_adapter.clk = clk;
										assign dcache_adapter.reset = reset;
										genvar _gv_j_15;
										for (_gv_j_15 = 0; _gv_j_15 < VX_gpu_pkg_DCACHE_CHANNELS; _gv_j_15 = _gv_j_15 + 1) begin : g_dcache_bus_if
											localparam j = _gv_j_15;
											// Trace: src/VX_mem_unit.sv:169:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((i * VX_gpu_pkg_DCACHE_CHANNELS) + j) + _mbase_dcache_bus_if].req_valid = dcache_bus_tmp_if[j].req_valid;
											// Trace: src/VX_mem_unit.sv:170:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((i * VX_gpu_pkg_DCACHE_CHANNELS) + j) + _mbase_dcache_bus_if].req_data = dcache_bus_tmp_if[j].req_data;
											// Trace: src/VX_mem_unit.sv:171:5
											assign dcache_bus_tmp_if[j].req_ready = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((i * VX_gpu_pkg_DCACHE_CHANNELS) + j) + _mbase_dcache_bus_if].req_ready;
											// Trace: src/VX_mem_unit.sv:172:5
											assign dcache_bus_tmp_if[j].rsp_valid = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((i * VX_gpu_pkg_DCACHE_CHANNELS) + j) + _mbase_dcache_bus_if].rsp_valid;
											// Trace: src/VX_mem_unit.sv:173:5
											assign dcache_bus_tmp_if[j].rsp_data = Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((i * VX_gpu_pkg_DCACHE_CHANNELS) + j) + _mbase_dcache_bus_if].rsp_data;
											// Trace: src/VX_mem_unit.sv:174:5
											assign Vortex.g_clusters[_gv_cluster_id_1].cluster.g_sockets[_gv_socket_id_1].socket.per_core_dcache_bus_if[((i * VX_gpu_pkg_DCACHE_CHANNELS) + j) + _mbase_dcache_bus_if].rsp_ready = dcache_bus_tmp_if[j].rsp_ready;
										end
									end
								end
								assign mem_unit.clk = clk;
								assign mem_unit.reset = reset;
							end
							assign core.clk = clk;
							assign core.reset = core_reset;
							assign per_core_busy[core_id] = core.busy;
						end
						// Trace: src/VX_socket.sv:316:5
						VX_pipe_register #(
							.DATAW(1),
							.RESETW(1),
							.DEPTH(1'd0)
						) __buffer_ex253(
							.clk(clk),
							.reset(reset),
							.enable(1'b1),
							.data_in(|per_core_busy),
							.data_out(busy)
						);
					end
					assign socket.clk = clk;
					assign socket.reset = socket_reset;
					assign per_socket_busy[socket_id] = socket.busy;
				end
				// Trace: src/VX_cluster.sv:86:5
				VX_pipe_register #(
					.DATAW(1),
					.RESETW(1),
					.DEPTH(1'd0)
				) __buffer_ex156(
					.clk(clk),
					.reset(reset),
					.enable(1'b1),
					.data_in(|per_socket_busy),
					.data_out(busy)
				);
			end
			assign cluster.clk = clk;
			assign cluster.reset = cluster_reset;
			assign per_cluster_busy[cluster_id] = cluster.busy;
		end
	endgenerate
	// Trace: src/Vortex.sv:115:5
	VX_pipe_register #(
		.DATAW(1),
		.RESETW(1),
		.DEPTH(1'd0)
	) __buffer_ex161(
		.clk(clk),
		.reset(reset),
		.enable(1'b1),
		.data_in(|per_cluster_busy),
		.data_out(busy)
	);
	// Trace: src/Vortex.sv:126:5
endmodule
module VX_scan (
	data_in,
	data_out
);
	// Trace: src/VX_scan.sv:2:15
	parameter N = 1;
	// Trace: src/VX_scan.sv:3:15
	parameter OP = "^";
	// Trace: src/VX_scan.sv:4:15
	parameter REVERSE = 0;
	// Trace: src/VX_scan.sv:6:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_scan.sv:7:5
	output wire [N - 1:0] data_out;
	// Trace: src/VX_scan.sv:9:5
	localparam LOGN = $clog2(N);
	// Trace: src/VX_scan.sv:10:5
	wire [(LOGN >= 0 ? ((LOGN + 1) * N) - 1 : ((1 - LOGN) * N) + ((LOGN * N) - 1)):(LOGN >= 0 ? 0 : LOGN * N)] t;
	// Trace: src/VX_scan.sv:11:5
	generate
		if (REVERSE != 0) begin : g_data_in_reverse
			// Trace: src/VX_scan.sv:12:9
			assign t[(LOGN >= 0 ? 0 : LOGN) * N+:N] = data_in;
		end
		else begin : g_data_in_no_reverse
			// Trace: src/VX_scan.sv:14:9
			function automatic [N - 1:0] _sv2v_strm_F2A76;
				input reg [(0 + N) - 1:0] inp;
				reg [(0 + N) - 1:0] _sv2v_strm_55E18_inp;
				reg [(0 + N) - 1:0] _sv2v_strm_55E18_out;
				integer _sv2v_strm_55E18_idx;
				begin
					_sv2v_strm_55E18_inp = {inp};
					for (_sv2v_strm_55E18_idx = 0; _sv2v_strm_55E18_idx <= ((0 + N) - 1); _sv2v_strm_55E18_idx = _sv2v_strm_55E18_idx + 1)
						_sv2v_strm_55E18_out[((0 + N) - 1) - _sv2v_strm_55E18_idx-:1] = _sv2v_strm_55E18_inp[_sv2v_strm_55E18_idx+:1];
					_sv2v_strm_F2A76 = ((0 + N) <= N ? _sv2v_strm_55E18_out << (N - (0 + N)) : _sv2v_strm_55E18_out >> ((0 + N) - N));
				end
			endfunction
			assign t[(LOGN >= 0 ? 0 : LOGN) * N+:N] = _sv2v_strm_F2A76({data_in});
		end
	endgenerate
	// Trace: src/VX_scan.sv:16:5
	function automatic [N - 1:0] sv2v_cast_AC047;
		input reg [N - 1:0] inp;
		sv2v_cast_AC047 = inp;
	endfunction
	generate
		if ((N == 2) && (OP == "&")) begin : g_scan_n2_and
			// Trace: src/VX_scan.sv:17:6
			assign t[(LOGN >= 0 ? LOGN : LOGN - LOGN) * N+:N] = {t[((LOGN >= 0 ? 0 : LOGN) * N) + 1], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 1-:2]};
		end
		else if ((N == 3) && (OP == "&")) begin : g_scan_n3_and
			// Trace: src/VX_scan.sv:19:6
			assign t[(LOGN >= 0 ? LOGN : LOGN - LOGN) * N+:N] = {t[((LOGN >= 0 ? 0 : LOGN) * N) + 2], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 2-:2], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 2-:3]};
		end
		else if ((N == 4) && (OP == "&")) begin : g_scan_n4_and
			// Trace: src/VX_scan.sv:21:6
			assign t[(LOGN >= 0 ? LOGN : LOGN - LOGN) * N+:N] = {t[((LOGN >= 0 ? 0 : LOGN) * N) + 3], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 3-:2], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 3-:3], &t[((LOGN >= 0 ? 0 : LOGN) * N) + 3-:4]};
		end
		else begin : g_scan
			// Trace: src/VX_scan.sv:23:9
			wire [N - 1:0] fill;
			genvar _gv_i_96;
			for (_gv_i_96 = 0; _gv_i_96 < LOGN; _gv_i_96 = _gv_i_96 + 1) begin : g_i
				localparam i = _gv_i_96;
				// Trace: src/VX_scan.sv:25:13
				wire [N - 1:0] shifted = sv2v_cast_AC047({fill, t[(LOGN >= 0 ? i : LOGN - i) * N+:N]} >> (1 << i));
				if (OP == "^") begin : g_xor
					// Trace: src/VX_scan.sv:27:11
					assign fill = {N {1'b0}};
					// Trace: src/VX_scan.sv:28:11
					assign t[(LOGN >= 0 ? i + 1 : LOGN - (i + 1)) * N+:N] = t[(LOGN >= 0 ? i : LOGN - i) * N+:N] ^ shifted;
				end
				else if (OP == "&") begin : g_and
					// Trace: src/VX_scan.sv:30:11
					assign fill = {N {1'b1}};
					// Trace: src/VX_scan.sv:31:11
					assign t[(LOGN >= 0 ? i + 1 : LOGN - (i + 1)) * N+:N] = t[(LOGN >= 0 ? i : LOGN - i) * N+:N] & shifted;
				end
				else if (OP == "|") begin : g_or
					// Trace: src/VX_scan.sv:33:11
					assign fill = {N {1'b0}};
					// Trace: src/VX_scan.sv:34:11
					assign t[(LOGN >= 0 ? i + 1 : LOGN - (i + 1)) * N+:N] = t[(LOGN >= 0 ? i : LOGN - i) * N+:N] | shifted;
				end
			end
		end
	endgenerate
	// Trace: src/VX_scan.sv:38:5
	generate
		if (REVERSE != 0) begin : g_data_out_reverse
			// Trace: src/VX_scan.sv:39:9
			assign data_out = t[(LOGN >= 0 ? LOGN : LOGN - LOGN) * N+:N];
		end
		else begin : g_data_out
			genvar _gv_i_97;
			for (_gv_i_97 = 0; _gv_i_97 < N; _gv_i_97 = _gv_i_97 + 1) begin : g_i
				localparam i = _gv_i_97;
				// Trace: src/VX_scan.sv:42:13
				assign data_out[i] = t[((LOGN >= 0 ? LOGN : LOGN - LOGN) * N) + ((N - 1) - i)];
			end
		end
	endgenerate
endmodule
module VX_stream_xbar (
	clk,
	reset,
	valid_in,
	data_in,
	sel_in,
	ready_in,
	valid_out,
	data_out,
	sel_out,
	ready_out,
	collisions
);
	// Trace: src/VX_stream_xbar.sv:2:15
	parameter NUM_INPUTS = 4;
	// Trace: src/VX_stream_xbar.sv:3:15
	parameter NUM_OUTPUTS = 4;
	// Trace: src/VX_stream_xbar.sv:4:15
	parameter DATAW = 4;
	// Trace: src/VX_stream_xbar.sv:5:15
	parameter ARBITER = "R";
	// Trace: src/VX_stream_xbar.sv:6:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_stream_xbar.sv:7:15
	parameter MAX_FANOUT = 8;
	// Trace: src/VX_stream_xbar.sv:8:15
	parameter PERF_CTR_BITS = $clog2(NUM_INPUTS + 1);
	// Trace: src/VX_stream_xbar.sv:9:15
	parameter IN_WIDTH = (NUM_INPUTS > 1 ? $clog2(NUM_INPUTS) : 1);
	// Trace: src/VX_stream_xbar.sv:10:15
	parameter OUT_WIDTH = (NUM_OUTPUTS > 1 ? $clog2(NUM_OUTPUTS) : 1);
	// Trace: src/VX_stream_xbar.sv:12:5
	input wire clk;
	// Trace: src/VX_stream_xbar.sv:13:5
	input wire reset;
	// Trace: src/VX_stream_xbar.sv:14:5
	input wire [NUM_INPUTS - 1:0] valid_in;
	// Trace: src/VX_stream_xbar.sv:15:5
	input wire [(NUM_INPUTS * DATAW) - 1:0] data_in;
	// Trace: src/VX_stream_xbar.sv:16:5
	input wire [(NUM_INPUTS * OUT_WIDTH) - 1:0] sel_in;
	// Trace: src/VX_stream_xbar.sv:17:5
	output wire [NUM_INPUTS - 1:0] ready_in;
	// Trace: src/VX_stream_xbar.sv:18:5
	output wire [NUM_OUTPUTS - 1:0] valid_out;
	// Trace: src/VX_stream_xbar.sv:19:5
	output wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out;
	// Trace: src/VX_stream_xbar.sv:20:5
	output wire [(NUM_OUTPUTS * IN_WIDTH) - 1:0] sel_out;
	// Trace: src/VX_stream_xbar.sv:21:5
	input wire [NUM_OUTPUTS - 1:0] ready_out;
	// Trace: src/VX_stream_xbar.sv:22:5
	output wire [PERF_CTR_BITS - 1:0] collisions;
	// Trace: src/VX_stream_xbar.sv:24:5
	generate
		if (NUM_INPUTS != 1) begin : g_multi_inputs
			if (NUM_OUTPUTS != 1) begin : g_multiple_outputs
				// Trace: src/VX_stream_xbar.sv:26:13
				wire [(NUM_INPUTS * NUM_OUTPUTS) - 1:0] per_output_valid_in;
				// Trace: src/VX_stream_xbar.sv:27:13
				wire [(NUM_OUTPUTS * NUM_INPUTS) - 1:0] per_output_valid_in_w;
				// Trace: src/VX_stream_xbar.sv:28:13
				wire [(NUM_OUTPUTS * NUM_INPUTS) - 1:0] per_output_ready_in;
				// Trace: src/VX_stream_xbar.sv:29:13
				wire [(NUM_INPUTS * NUM_OUTPUTS) - 1:0] per_output_ready_in_w;
				// Trace: src/VX_stream_xbar.sv:30:13
				VX_transpose #(
					.N(NUM_OUTPUTS),
					.M(NUM_INPUTS)
				) rdy_in_transpose(
					.data_in(per_output_ready_in),
					.data_out(per_output_ready_in_w)
				);
				genvar _gv_i_105;
				for (_gv_i_105 = 0; _gv_i_105 < NUM_INPUTS; _gv_i_105 = _gv_i_105 + 1) begin : g_ready_in
					localparam i = _gv_i_105;
					// Trace: src/VX_stream_xbar.sv:38:17
					assign ready_in[i] = |per_output_ready_in_w[i * NUM_OUTPUTS+:NUM_OUTPUTS];
				end
				genvar _gv_i_106;
				for (_gv_i_106 = 0; _gv_i_106 < NUM_INPUTS; _gv_i_106 = _gv_i_106 + 1) begin : g_sel_in_demux
					localparam i = _gv_i_106;
					// Trace: src/VX_stream_xbar.sv:41:17
					VX_demux #(
						.DATAW(1),
						.N(NUM_OUTPUTS)
					) sel_in_demux(
						.sel_in(sel_in[i * OUT_WIDTH+:OUT_WIDTH]),
						.data_in(valid_in[i]),
						.data_out(per_output_valid_in[i * NUM_OUTPUTS+:NUM_OUTPUTS])
					);
				end
				// Trace: src/VX_stream_xbar.sv:50:13
				VX_transpose #(
					.N(NUM_INPUTS),
					.M(NUM_OUTPUTS)
				) val_in_transpose(
					.data_in(per_output_valid_in),
					.data_out(per_output_valid_in_w)
				);
				genvar _gv_i_107;
				for (_gv_i_107 = 0; _gv_i_107 < NUM_OUTPUTS; _gv_i_107 = _gv_i_107 + 1) begin : g_xbar_arbs
					localparam i = _gv_i_107;
					// Trace: src/VX_stream_xbar.sv:58:17
					VX_stream_arb #(
						.NUM_INPUTS(NUM_INPUTS),
						.NUM_OUTPUTS(1),
						.DATAW(DATAW),
						.ARBITER(ARBITER),
						.MAX_FANOUT(MAX_FANOUT),
						.OUT_BUF(OUT_BUF)
					) xbar_arb(
						.clk(clk),
						.reset(reset),
						.valid_in(per_output_valid_in_w[i * NUM_INPUTS+:NUM_INPUTS]),
						.data_in(data_in),
						.ready_in(per_output_ready_in[i * NUM_INPUTS+:NUM_INPUTS]),
						.valid_out(valid_out[i]),
						.data_out(data_out[i * DATAW+:DATAW]),
						.sel_out(sel_out[i * IN_WIDTH+:IN_WIDTH]),
						.ready_out(ready_out[i])
					);
				end
			end
			else begin : g_one_output
				// Trace: src/VX_stream_xbar.sv:78:13
				VX_stream_arb #(
					.NUM_INPUTS(NUM_INPUTS),
					.NUM_OUTPUTS(1),
					.DATAW(DATAW),
					.ARBITER(ARBITER),
					.MAX_FANOUT(MAX_FANOUT),
					.OUT_BUF(OUT_BUF)
				) xbar_arb(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_in),
					.data_in(data_in),
					.ready_in(ready_in),
					.valid_out(valid_out),
					.data_out(data_out),
					.sel_out(sel_out),
					.ready_out(ready_out)
				);
			end
		end
		else if (NUM_OUTPUTS != 1) begin : g_single_input
			// Trace: src/VX_stream_xbar.sv:98:9
			wire [NUM_OUTPUTS - 1:0] valid_out_w;
			wire [NUM_OUTPUTS - 1:0] ready_out_w;
			// Trace: src/VX_stream_xbar.sv:99:9
			wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out_w;
			// Trace: src/VX_stream_xbar.sv:100:9
			VX_demux #(
				.DATAW(1),
				.N(NUM_OUTPUTS)
			) sel_in_demux(
				.sel_in(sel_in[0+:OUT_WIDTH]),
				.data_in(valid_in[0]),
				.data_out(valid_out_w)
			);
			// Trace: src/VX_stream_xbar.sv:108:9
			assign ready_in[0] = ready_out_w[sel_in[0+:OUT_WIDTH]];
			// Trace: src/VX_stream_xbar.sv:109:9
			assign data_out_w = {NUM_OUTPUTS {data_in[0+:DATAW]}};
			genvar _gv_i_108;
			for (_gv_i_108 = 0; _gv_i_108 < NUM_OUTPUTS; _gv_i_108 = _gv_i_108 + 1) begin : g_out_buf
				localparam i = _gv_i_108;
				// Trace: src/VX_stream_xbar.sv:111:13
				VX_elastic_buffer #(
					.DATAW(DATAW),
					.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
					.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2)),
					.LUTRAM((OUT_BUF & 8) != 0)
				) out_buf(
					.clk(clk),
					.reset(reset),
					.valid_in(valid_out_w[i]),
					.ready_in(ready_out_w[i]),
					.data_in(data_out_w[i * DATAW+:DATAW]),
					.data_out(data_out[i * DATAW+:DATAW]),
					.valid_out(valid_out[i]),
					.ready_out(ready_out[i])
				);
			end
			// Trace: src/VX_stream_xbar.sv:127:9
			assign sel_out = 0;
		end
		else begin : g_passthru
			// Trace: src/VX_stream_xbar.sv:129:9
			VX_elastic_buffer #(
				.DATAW(DATAW),
				.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
				.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2)),
				.LUTRAM((OUT_BUF & 8) != 0)
			) out_buf(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_in),
				.ready_in(ready_in),
				.data_in(data_in),
				.data_out(data_out),
				.valid_out(valid_out),
				.ready_out(ready_out)
			);
			// Trace: src/VX_stream_xbar.sv:144:9
			assign sel_out = 0;
		end
	endgenerate
	// Trace: src/VX_stream_xbar.sv:146:5
	reg [NUM_INPUTS - 1:0] per_cycle_collision;
	reg [NUM_INPUTS - 1:0] per_cycle_collision_r;
	// Trace: src/VX_stream_xbar.sv:147:5
	wire [$clog2(NUM_INPUTS + 1) - 1:0] collision_count;
	// Trace: src/VX_stream_xbar.sv:148:5
	reg [PERF_CTR_BITS - 1:0] collisions_r;
	// Trace: src/VX_stream_xbar.sv:149:5
	always @(*) begin
		// Trace: src/VX_stream_xbar.sv:150:9
		per_cycle_collision = 1'sb0;
		// Trace: src/VX_stream_xbar.sv:151:9
		begin : sv2v_autoblock_1
			// Trace: src/VX_stream_xbar.sv:151:14
			integer i;
			// Trace: src/VX_stream_xbar.sv:151:14
			for (i = 0; i < NUM_INPUTS; i = i + 1)
				begin
					// Trace: src/VX_stream_xbar.sv:152:13
					begin : sv2v_autoblock_2
						// Trace: src/VX_stream_xbar.sv:152:18
						integer j;
						// Trace: src/VX_stream_xbar.sv:152:18
						for (j = i + 1; j < NUM_INPUTS; j = j + 1)
							begin
								// Trace: src/VX_stream_xbar.sv:153:17
								per_cycle_collision[i] = per_cycle_collision[i] | (((valid_in[i] && valid_in[j]) && (sel_in[i * OUT_WIDTH+:OUT_WIDTH] == sel_in[j * OUT_WIDTH+:OUT_WIDTH])) && (ready_in[i] | ready_in[j]));
							end
					end
				end
		end
	end
	// Trace: src/VX_stream_xbar.sv:160:5
	// rewrote reg-to-output bindings
	wire [NUM_INPUTS:1] sv2v_tmp___buffer_ex220_data_out;
	always @(*) per_cycle_collision_r = sv2v_tmp___buffer_ex220_data_out;
	VX_pipe_register #(
		.DATAW(NUM_INPUTS),
		.RESETW(NUM_INPUTS),
		.DEPTH(1)
	) __buffer_ex220(
		.clk(clk),
		.reset(reset),
		.enable(1'b1),
		.data_in(per_cycle_collision),
		.data_out(sv2v_tmp___buffer_ex220_data_out)
	);
	// Trace: src/VX_stream_xbar.sv:171:5
	VX_popcount #(
		.N(NUM_INPUTS),
		.MODEL(1)
	) __pop_count_ex221(
		.data_in(per_cycle_collision_r),
		.data_out(collision_count)
	);
	// Trace: src/VX_stream_xbar.sv:178:5
	function automatic [PERF_CTR_BITS - 1:0] sv2v_cast_8BEE5;
		input reg [PERF_CTR_BITS - 1:0] inp;
		sv2v_cast_8BEE5 = inp;
	endfunction
	always @(posedge clk)
		// Trace: src/VX_stream_xbar.sv:179:9
		if (reset)
			// Trace: src/VX_stream_xbar.sv:180:13
			collisions_r <= 1'sb0;
		else
			// Trace: src/VX_stream_xbar.sv:182:13
			collisions_r <= collisions_r + sv2v_cast_8BEE5(collision_count);
	// Trace: src/VX_stream_xbar.sv:185:5
	assign collisions = collisions_r;
endmodule
// removed interface: VX_schedule_if
// removed module with interface ports: VX_mem_switch
// removed module with interface ports: VX_lsu_slice
module VX_stream_omega (
	clk,
	reset,
	valid_in,
	data_in,
	sel_in,
	ready_in,
	valid_out,
	data_out,
	sel_out,
	ready_out,
	collisions
);
	// Trace: src/VX_stream_omega.sv:2:15
	parameter NUM_INPUTS = 4;
	// Trace: src/VX_stream_omega.sv:3:15
	parameter NUM_OUTPUTS = 4;
	// Trace: src/VX_stream_omega.sv:4:15
	parameter RADIX = 2;
	// Trace: src/VX_stream_omega.sv:5:15
	parameter DATAW = 4;
	// Trace: src/VX_stream_omega.sv:6:15
	parameter ARBITER = "R";
	// Trace: src/VX_stream_omega.sv:7:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_stream_omega.sv:8:15
	parameter MAX_FANOUT = 8;
	// Trace: src/VX_stream_omega.sv:9:15
	parameter PERF_CTR_BITS = 32;
	// Trace: src/VX_stream_omega.sv:10:15
	parameter IN_WIDTH = (NUM_INPUTS > 1 ? $clog2(NUM_INPUTS) : 1);
	// Trace: src/VX_stream_omega.sv:11:15
	parameter OUT_WIDTH = (NUM_OUTPUTS > 1 ? $clog2(NUM_OUTPUTS) : 1);
	// Trace: src/VX_stream_omega.sv:13:5
	input wire clk;
	// Trace: src/VX_stream_omega.sv:14:5
	input wire reset;
	// Trace: src/VX_stream_omega.sv:15:5
	input wire [NUM_INPUTS - 1:0] valid_in;
	// Trace: src/VX_stream_omega.sv:16:5
	input wire [(NUM_INPUTS * DATAW) - 1:0] data_in;
	// Trace: src/VX_stream_omega.sv:17:5
	input wire [(NUM_INPUTS * OUT_WIDTH) - 1:0] sel_in;
	// Trace: src/VX_stream_omega.sv:18:5
	output wire [NUM_INPUTS - 1:0] ready_in;
	// Trace: src/VX_stream_omega.sv:19:5
	output wire [NUM_OUTPUTS - 1:0] valid_out;
	// Trace: src/VX_stream_omega.sv:20:5
	output wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out;
	// Trace: src/VX_stream_omega.sv:21:5
	output wire [(NUM_OUTPUTS * IN_WIDTH) - 1:0] sel_out;
	// Trace: src/VX_stream_omega.sv:22:5
	input wire [NUM_OUTPUTS - 1:0] ready_out;
	// Trace: src/VX_stream_omega.sv:23:5
	output wire [PERF_CTR_BITS - 1:0] collisions;
	// Trace: src/VX_stream_omega.sv:25:5
	function automatic [DATAW - 1:0] sv2v_cast_8E21C;
		input reg [DATAW - 1:0] inp;
		sv2v_cast_8E21C = inp;
	endfunction
	function automatic signed [IN_WIDTH - 1:0] sv2v_cast_314B8_signed;
		input reg signed [IN_WIDTH - 1:0] inp;
		sv2v_cast_314B8_signed = inp;
	endfunction
	function automatic [IN_WIDTH - 1:0] sv2v_cast_314B8;
		input reg [IN_WIDTH - 1:0] inp;
		sv2v_cast_314B8 = inp;
	endfunction
	function automatic [PERF_CTR_BITS - 1:0] sv2v_cast_8BEE5;
		input reg [PERF_CTR_BITS - 1:0] inp;
		sv2v_cast_8BEE5 = inp;
	endfunction
	generate
		if ((NUM_INPUTS <= RADIX) && (NUM_OUTPUTS <= RADIX)) begin : g_fallback
			// Trace: src/VX_stream_omega.sv:26:9
			VX_stream_xbar #(
				.NUM_INPUTS(NUM_INPUTS),
				.NUM_OUTPUTS(NUM_OUTPUTS),
				.DATAW(DATAW),
				.ARBITER(ARBITER),
				.OUT_BUF(OUT_BUF),
				.MAX_FANOUT(MAX_FANOUT),
				.PERF_CTR_BITS(PERF_CTR_BITS)
			) xbar_switch(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_in),
				.data_in(data_in),
				.sel_in(sel_in),
				.ready_in(ready_in),
				.valid_out(valid_out),
				.data_out(data_out),
				.sel_out(sel_out),
				.ready_out(ready_out),
				.collisions(collisions)
			);
		end
		else begin : g_omega
			// Trace: src/VX_stream_omega.sv:48:9
			localparam RADIX_LG = (RADIX > 1 ? $clog2(RADIX) : 1);
			// Trace: src/VX_stream_omega.sv:49:9
			localparam N_INPUTS_M = (NUM_INPUTS > NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
			// Trace: src/VX_stream_omega.sv:50:9
			localparam N_INPUTS_LG = (($clog2(N_INPUTS_M) + RADIX_LG) - 1) / RADIX_LG;
			// Trace: src/VX_stream_omega.sv:51:9
			localparam N_INPUTS = RADIX ** N_INPUTS_LG;
			// Trace: src/VX_stream_omega.sv:52:9
			localparam NUM_STAGES = (N_INPUTS > 1 ? $clog2(N_INPUTS) : 1) / RADIX_LG;
			// Trace: src/VX_stream_omega.sv:53:9
			localparam NUM_SWITCHES = N_INPUTS / RADIX;
			// Trace: src/VX_stream_omega.sv:54:9
			// removed localparam type omega_t
			// Trace: src/VX_stream_omega.sv:59:9
			wire [((NUM_STAGES * NUM_SWITCHES) * RADIX) - 1:0] switch_valid_in;
			wire [((NUM_STAGES * NUM_SWITCHES) * RADIX) - 1:0] switch_valid_out;
			// Trace: src/VX_stream_omega.sv:60:9
			wire [(((NUM_STAGES * NUM_SWITCHES) * RADIX) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)) - 1:0] switch_data_in;
			wire [(((NUM_STAGES * NUM_SWITCHES) * RADIX) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)) - 1:0] switch_data_out;
			// Trace: src/VX_stream_omega.sv:61:9
			wire [(((NUM_STAGES * NUM_SWITCHES) * RADIX) * RADIX_LG) - 1:0] switch_sel_in;
			// Trace: src/VX_stream_omega.sv:62:9
			wire [((NUM_STAGES * NUM_SWITCHES) * RADIX) - 1:0] switch_ready_in;
			wire [((NUM_STAGES * NUM_SWITCHES) * RADIX) - 1:0] switch_ready_out;
			genvar _gv_i_120;
			for (_gv_i_120 = 0; _gv_i_120 < N_INPUTS; _gv_i_120 = _gv_i_120 + 1) begin : g_tie_inputs
				localparam i = _gv_i_120;
				// Trace: src/VX_stream_omega.sv:64:13
				localparam DST_IDX = ((i << 1) | (i >> (N_INPUTS_LG - 1))) & (N_INPUTS - 1);
				// Trace: src/VX_stream_omega.sv:65:13
				localparam switch = DST_IDX / RADIX;
				// Trace: src/VX_stream_omega.sv:66:13
				localparam port = DST_IDX % RADIX;
				if (i < NUM_INPUTS) begin : g_valid
					// Trace: src/VX_stream_omega.sv:68:17
					assign switch_valid_in[((0 + switch) * RADIX) + port] = valid_in[i];
					// Trace: src/VX_stream_omega.sv:69:17
					function automatic [N_INPUTS_LG - 1:0] sv2v_cast_51E45;
						input reg [N_INPUTS_LG - 1:0] inp;
						sv2v_cast_51E45 = inp;
					endfunction
					function automatic [N_INPUTS_LG - 1:0] sv2v_cast_43513;
						input reg [N_INPUTS_LG - 1:0] inp;
						sv2v_cast_43513 = inp;
					endfunction
					assign switch_data_in[(((0 + switch) * RADIX) + port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)+:(N_INPUTS_LG + DATAW) + IN_WIDTH] = {sv2v_cast_43513(sv2v_cast_51E45(sel_in[i * OUT_WIDTH+:OUT_WIDTH])), sv2v_cast_8E21C(data_in[i * DATAW+:DATAW]), sv2v_cast_314B8(sv2v_cast_314B8_signed(i))};
					// Trace: src/VX_stream_omega.sv:74:17
					assign ready_in[i] = switch_ready_in[((0 + switch) * RADIX) + port];
				end
				else begin : g_padding
					// Trace: src/VX_stream_omega.sv:76:17
					assign switch_valid_in[((0 + switch) * RADIX) + port] = 0;
					// Trace: src/VX_stream_omega.sv:77:17
					assign switch_data_in[(((0 + switch) * RADIX) + port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)+:(N_INPUTS_LG + DATAW) + IN_WIDTH] = 1'sbx;
				end
			end
			genvar _gv_stage_1;
			for (_gv_stage_1 = 0; _gv_stage_1 < NUM_STAGES; _gv_stage_1 = _gv_stage_1 + 1) begin : g_sel_in
				localparam stage = _gv_stage_1;
				genvar _gv_switch_1;
				for (_gv_switch_1 = 0; _gv_switch_1 < NUM_SWITCHES; _gv_switch_1 = _gv_switch_1 + 1) begin : g_switches
					localparam switch = _gv_switch_1;
					genvar _gv_port_1;
					for (_gv_port_1 = 0; _gv_port_1 < RADIX; _gv_port_1 = _gv_port_1 + 1) begin : g_ports
						localparam port = _gv_port_1;
						// Trace: src/VX_stream_omega.sv:83:21
						assign switch_sel_in[((((stage * NUM_SWITCHES) + switch) * RADIX) + port) * RADIX_LG+:RADIX_LG] = switch_data_in[(((((stage * NUM_SWITCHES) + switch) * RADIX) + port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)) + ((N_INPUTS_LG + (DATAW + (IN_WIDTH - 1))) - ((N_INPUTS_LG - 1) - (((NUM_STAGES - 1) - stage) * RADIX_LG)))+:RADIX_LG];
					end
				end
			end
			genvar _gv_stage_2;
			for (_gv_stage_2 = 0; _gv_stage_2 < (NUM_STAGES - 1); _gv_stage_2 = _gv_stage_2 + 1) begin : g_stages
				localparam stage = _gv_stage_2;
				genvar _gv_switch_2;
				for (_gv_switch_2 = 0; _gv_switch_2 < NUM_SWITCHES; _gv_switch_2 = _gv_switch_2 + 1) begin : g_switches
					localparam switch = _gv_switch_2;
					genvar _gv_port_2;
					for (_gv_port_2 = 0; _gv_port_2 < RADIX; _gv_port_2 = _gv_port_2 + 1) begin : g_ports
						localparam port = _gv_port_2;
						// Trace: src/VX_stream_omega.sv:90:21
						localparam lane = (switch * RADIX) + port;
						// Trace: src/VX_stream_omega.sv:91:21
						localparam dst_lane = ((lane << 1) | (lane >> (N_INPUTS_LG - 1))) & (N_INPUTS - 1);
						// Trace: src/VX_stream_omega.sv:92:21
						localparam dst_switch = dst_lane / RADIX;
						// Trace: src/VX_stream_omega.sv:93:21
						localparam dst_port = dst_lane % RADIX;
						// Trace: src/VX_stream_omega.sv:94:21
						assign switch_valid_in[((((stage + 1) * NUM_SWITCHES) + dst_switch) * RADIX) + dst_port] = switch_valid_out[(((stage * NUM_SWITCHES) + switch) * RADIX) + port];
						// Trace: src/VX_stream_omega.sv:95:21
						assign switch_data_in[(((((stage + 1) * NUM_SWITCHES) + dst_switch) * RADIX) + dst_port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)+:(N_INPUTS_LG + DATAW) + IN_WIDTH] = switch_data_out[((((stage * NUM_SWITCHES) + switch) * RADIX) + port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)+:(N_INPUTS_LG + DATAW) + IN_WIDTH];
						// Trace: src/VX_stream_omega.sv:96:21
						assign switch_ready_out[(((stage * NUM_SWITCHES) + switch) * RADIX) + port] = switch_ready_in[((((stage + 1) * NUM_SWITCHES) + dst_switch) * RADIX) + dst_port];
					end
				end
			end
			genvar _gv_switch_3;
			for (_gv_switch_3 = 0; _gv_switch_3 < NUM_SWITCHES; _gv_switch_3 = _gv_switch_3 + 1) begin : g_switches
				localparam switch = _gv_switch_3;
				genvar _gv_stage_3;
				for (_gv_stage_3 = 0; _gv_stage_3 < NUM_STAGES; _gv_stage_3 = _gv_stage_3 + 1) begin : g_stages
					localparam stage = _gv_stage_3;
					// Trace: src/VX_stream_omega.sv:102:17
					VX_stream_xbar #(
						.NUM_INPUTS(RADIX),
						.NUM_OUTPUTS(RADIX),
						.DATAW((N_INPUTS_LG + DATAW) + IN_WIDTH),
						.ARBITER(ARBITER),
						.OUT_BUF(OUT_BUF),
						.MAX_FANOUT(MAX_FANOUT),
						.PERF_CTR_BITS(PERF_CTR_BITS)
					) xbar_switch(
						.clk(clk),
						.reset(reset),
						.valid_in(switch_valid_in[((stage * NUM_SWITCHES) + switch) * RADIX+:RADIX]),
						.data_in(switch_data_in[((N_INPUTS_LG + DATAW) + IN_WIDTH) * (((stage * NUM_SWITCHES) + switch) * RADIX)+:((N_INPUTS_LG + DATAW) + IN_WIDTH) * RADIX]),
						.sel_in(switch_sel_in[RADIX_LG * (((stage * NUM_SWITCHES) + switch) * RADIX)+:RADIX_LG * RADIX]),
						.ready_in(switch_ready_in[((stage * NUM_SWITCHES) + switch) * RADIX+:RADIX]),
						.valid_out(switch_valid_out[((stage * NUM_SWITCHES) + switch) * RADIX+:RADIX]),
						.data_out(switch_data_out[((N_INPUTS_LG + DATAW) + IN_WIDTH) * (((stage * NUM_SWITCHES) + switch) * RADIX)+:((N_INPUTS_LG + DATAW) + IN_WIDTH) * RADIX]),
						.sel_out(),
						.ready_out(switch_ready_out[((stage * NUM_SWITCHES) + switch) * RADIX+:RADIX]),
						.collisions()
					);
				end
			end
			genvar _gv_i_121;
			for (_gv_i_121 = 0; _gv_i_121 < N_INPUTS; _gv_i_121 = _gv_i_121 + 1) begin : g_tie_outputs
				localparam i = _gv_i_121;
				// Trace: src/VX_stream_omega.sv:126:13
				localparam switch = i / RADIX;
				// Trace: src/VX_stream_omega.sv:127:13
				localparam port = i % RADIX;
				if (i < NUM_OUTPUTS) begin : g_valid
					// Trace: src/VX_stream_omega.sv:129:17
					assign valid_out[i] = switch_valid_out[((((NUM_STAGES - 1) * NUM_SWITCHES) + switch) * RADIX) + port];
					// Trace: src/VX_stream_omega.sv:130:17
					assign data_out[i * DATAW+:DATAW] = switch_data_out[((((((NUM_STAGES - 1) * NUM_SWITCHES) + switch) * RADIX) + port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)) + (DATAW + (IN_WIDTH - 1))-:((DATAW + (IN_WIDTH - 1)) >= (IN_WIDTH + 0) ? ((DATAW + (IN_WIDTH - 1)) - (IN_WIDTH + 0)) + 1 : ((IN_WIDTH + 0) - (DATAW + (IN_WIDTH - 1))) + 1)];
					// Trace: src/VX_stream_omega.sv:131:17
					assign sel_out[i * IN_WIDTH+:IN_WIDTH] = switch_data_out[((((((NUM_STAGES - 1) * NUM_SWITCHES) + switch) * RADIX) + port) * ((N_INPUTS_LG + DATAW) + IN_WIDTH)) + (IN_WIDTH - 1)-:IN_WIDTH];
					// Trace: src/VX_stream_omega.sv:132:17
					assign switch_ready_out[((((NUM_STAGES - 1) * NUM_SWITCHES) + switch) * RADIX) + port] = ready_out[i];
				end
				else begin : g_padding
					// Trace: src/VX_stream_omega.sv:134:17
					assign switch_ready_out[((((NUM_STAGES - 1) * NUM_SWITCHES) + switch) * RADIX) + port] = 0;
				end
			end
			// Trace: src/VX_stream_omega.sv:137:9
			reg [((NUM_STAGES * NUM_SWITCHES) * RADIX) - 1:0] per_cycle_collision;
			reg [((NUM_STAGES * NUM_SWITCHES) * RADIX) - 1:0] per_cycle_collision_r;
			// Trace: src/VX_stream_omega.sv:138:9
			wire [$clog2(((NUM_STAGES * NUM_SWITCHES) * RADIX) + 1) - 1:0] collision_count;
			// Trace: src/VX_stream_omega.sv:139:9
			reg [PERF_CTR_BITS - 1:0] collisions_r;
			// Trace: src/VX_stream_omega.sv:140:9
			always @(*) begin
				// Trace: src/VX_stream_omega.sv:141:13
				per_cycle_collision = 0;
				// Trace: src/VX_stream_omega.sv:142:13
				begin : sv2v_autoblock_1
					// Trace: src/VX_stream_omega.sv:142:18
					integer stage;
					// Trace: src/VX_stream_omega.sv:142:18
					for (stage = 0; stage < NUM_STAGES; stage = stage + 1)
						begin
							// Trace: src/VX_stream_omega.sv:143:17
							begin : sv2v_autoblock_2
								// Trace: src/VX_stream_omega.sv:143:22
								integer switch;
								// Trace: src/VX_stream_omega.sv:143:22
								for (switch = 0; switch < NUM_SWITCHES; switch = switch + 1)
									begin
										// Trace: src/VX_stream_omega.sv:144:21
										begin : sv2v_autoblock_3
											// Trace: src/VX_stream_omega.sv:144:26
											integer port_a;
											// Trace: src/VX_stream_omega.sv:144:26
											for (port_a = 0; port_a < RADIX; port_a = port_a + 1)
												begin
													// Trace: src/VX_stream_omega.sv:145:25
													begin : sv2v_autoblock_4
														// Trace: src/VX_stream_omega.sv:145:30
														integer port_b;
														// Trace: src/VX_stream_omega.sv:145:30
														for (port_b = port_a + 1; port_b < RADIX; port_b = port_b + 1)
															begin
																// Trace: src/VX_stream_omega.sv:146:29
																per_cycle_collision[(((stage * NUM_SWITCHES) + switch) * RADIX) + port_a] = per_cycle_collision[(((stage * NUM_SWITCHES) + switch) * RADIX) + port_a] | (((switch_valid_in[(((stage * NUM_SWITCHES) + switch) * RADIX) + port_a] && switch_valid_in[(((stage * NUM_SWITCHES) + switch) * RADIX) + port_b]) && (switch_sel_in[((((stage * NUM_SWITCHES) + switch) * RADIX) + port_a) * RADIX_LG+:RADIX_LG] == switch_sel_in[((((stage * NUM_SWITCHES) + switch) * RADIX) + port_b) * RADIX_LG+:RADIX_LG])) && (switch_ready_in[(((stage * NUM_SWITCHES) + switch) * RADIX) + port_a] | switch_ready_in[(((stage * NUM_SWITCHES) + switch) * RADIX) + port_b]));
															end
													end
												end
										end
									end
							end
						end
				end
			end
			// Trace: src/VX_stream_omega.sv:155:5
			// rewrote reg-to-output bindings
			wire [(NUM_STAGES * NUM_SWITCHES) * RADIX:1] sv2v_tmp___buffer_ex200_data_out;
			always @(*) per_cycle_collision_r = sv2v_tmp___buffer_ex200_data_out;
			VX_pipe_register #(
				.DATAW((NUM_STAGES * NUM_SWITCHES) * RADIX),
				.RESETW((NUM_STAGES * NUM_SWITCHES) * RADIX),
				.DEPTH(1)
			) __buffer_ex200(
				.clk(clk),
				.reset(reset),
				.enable(1'b1),
				.data_in(per_cycle_collision),
				.data_out(sv2v_tmp___buffer_ex200_data_out)
			);
			// Trace: src/VX_stream_omega.sv:166:5
			VX_popcount #(
				.N((NUM_STAGES * NUM_SWITCHES) * RADIX),
				.MODEL(1)
			) __pop_count_ex201(
				.data_in(per_cycle_collision_r),
				.data_out(collision_count)
			);
			// Trace: src/VX_stream_omega.sv:173:9
			always @(posedge clk)
				// Trace: src/VX_stream_omega.sv:174:13
				if (reset)
					// Trace: src/VX_stream_omega.sv:175:17
					collisions_r <= 1'sb0;
				else
					// Trace: src/VX_stream_omega.sv:177:17
					collisions_r <= collisions_r + sv2v_cast_8BEE5(collision_count);
			// Trace: src/VX_stream_omega.sv:180:9
			assign collisions = collisions_r;
		end
	endgenerate
endmodule
// removed module with interface ports: VX_issue_slice
module VX_sp_ram (
	clk,
	reset,
	read,
	write,
	wren,
	addr,
	wdata,
	rdata
);
	// Trace: src/VX_sp_ram.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_sp_ram.sv:3:15
	parameter SIZE = 1;
	// Trace: src/VX_sp_ram.sv:4:15
	parameter WRENW = 1;
	// Trace: src/VX_sp_ram.sv:5:15
	parameter OUT_REG = 0;
	// Trace: src/VX_sp_ram.sv:6:15
	parameter LUTRAM = 0;
	// Trace: src/VX_sp_ram.sv:7:15
	parameter RDW_MODE = "W";
	// Trace: src/VX_sp_ram.sv:8:15
	parameter RADDR_REG = 0;
	// Trace: src/VX_sp_ram.sv:9:15
	parameter RADDR_RESET = 0;
	// Trace: src/VX_sp_ram.sv:10:15
	parameter RDW_ASSERT = 0;
	// Trace: src/VX_sp_ram.sv:11:15
	parameter RESET_RAM = 0;
	// Trace: src/VX_sp_ram.sv:12:15
	parameter INIT_ENABLE = 0;
	// Trace: src/VX_sp_ram.sv:13:15
	parameter INIT_FILE = "";
	// Trace: src/VX_sp_ram.sv:14:15
	parameter [DATAW - 1:0] INIT_VALUE = 0;
	// Trace: src/VX_sp_ram.sv:15:15
	parameter ADDRW = (SIZE > 1 ? $clog2(SIZE) : 1);
	// Trace: src/VX_sp_ram.sv:17:5
	input wire clk;
	// Trace: src/VX_sp_ram.sv:18:5
	input wire reset;
	// Trace: src/VX_sp_ram.sv:19:5
	input wire read;
	// Trace: src/VX_sp_ram.sv:20:5
	input wire write;
	// Trace: src/VX_sp_ram.sv:21:5
	input wire [WRENW - 1:0] wren;
	// Trace: src/VX_sp_ram.sv:22:5
	input wire [ADDRW - 1:0] addr;
	// Trace: src/VX_sp_ram.sv:23:5
	input wire [DATAW - 1:0] wdata;
	// Trace: src/VX_sp_ram.sv:24:5
	output wire [DATAW - 1:0] rdata;
	// Trace: src/VX_sp_ram.sv:26:5
	localparam WSELW = DATAW / WRENW;
	// Trace: src/VX_sp_ram.sv:27:5
	localparam FORCE_BRAM = !LUTRAM && ((((SIZE >= 64) || (DATAW >= 16)) || ((SIZE * DATAW) >= 512)) && ((SIZE * DATAW) >= 64));
	// Trace: src/VX_sp_ram.sv:28:5
	generate
		if (OUT_REG) begin : g_sync
			if (FORCE_BRAM) begin : g_bram
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:32:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:35:13
								initial begin
									// Trace: src/VX_sp_ram.sv:35:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:37:13
								initial begin
									// Trace: src/VX_sp_ram.sv:38:17
									begin : sv2v_autoblock_1
										// Trace: src/VX_sp_ram.sv:38:22
										integer i;
										// Trace: src/VX_sp_ram.sv:38:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:39:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:44:21
						reg [ADDRW - 1:0] addr_r;
						// Trace: src/VX_sp_ram.sv:45:21
						always @(posedge clk) begin
							// Trace: src/VX_sp_ram.sv:46:29
							if (write)
								// Trace: src/VX_sp_ram.sv:47:33
								begin : sv2v_autoblock_2
									// Trace: src/VX_sp_ram.sv:47:38
									integer i;
									// Trace: src/VX_sp_ram.sv:47:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:48:37
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:49:41
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							if (read)
								// Trace: src/VX_sp_ram.sv:54:29
								addr_r <= addr;
						end
						// Trace: src/VX_sp_ram.sv:57:21
						assign rdata = ram[addr_r];
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:59:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:62:13
								initial begin
									// Trace: src/VX_sp_ram.sv:62:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:64:13
								initial begin
									// Trace: src/VX_sp_ram.sv:65:17
									begin : sv2v_autoblock_3
										// Trace: src/VX_sp_ram.sv:65:22
										integer i;
										// Trace: src/VX_sp_ram.sv:65:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:66:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:71:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:72:21
						always @(posedge clk) begin
							// Trace: src/VX_sp_ram.sv:73:25
							if (write)
								// Trace: src/VX_sp_ram.sv:74:29
								ram[addr] <= wdata;
							if (read) begin
								begin
									// Trace: src/VX_sp_ram.sv:77:29
									if (write)
										// Trace: src/VX_sp_ram.sv:78:33
										rdata_r <= wdata;
									else
										// Trace: src/VX_sp_ram.sv:80:33
										rdata_r <= ram[addr];
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:84:21
						assign rdata = rdata_r;
					end
				end
				else if (RDW_MODE == "R") begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:88:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:91:13
								initial begin
									// Trace: src/VX_sp_ram.sv:91:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:93:13
								initial begin
									// Trace: src/VX_sp_ram.sv:94:17
									begin : sv2v_autoblock_4
										// Trace: src/VX_sp_ram.sv:94:22
										integer i;
										// Trace: src/VX_sp_ram.sv:94:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:95:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:100:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:101:21
						always @(posedge clk) begin
							// Trace: src/VX_sp_ram.sv:102:29
							if (write)
								// Trace: src/VX_sp_ram.sv:103:33
								begin : sv2v_autoblock_5
									// Trace: src/VX_sp_ram.sv:103:38
									integer i;
									// Trace: src/VX_sp_ram.sv:103:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:104:37
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:105:41
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							if (read)
								// Trace: src/VX_sp_ram.sv:110:29
								rdata_r <= ram[addr];
						end
						// Trace: src/VX_sp_ram.sv:113:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:115:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:118:13
								initial begin
									// Trace: src/VX_sp_ram.sv:118:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:120:13
								initial begin
									// Trace: src/VX_sp_ram.sv:121:17
									begin : sv2v_autoblock_6
										// Trace: src/VX_sp_ram.sv:121:22
										integer i;
										// Trace: src/VX_sp_ram.sv:121:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:122:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:127:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:128:21
						always @(posedge clk) begin
							// Trace: src/VX_sp_ram.sv:129:25
							if (write)
								// Trace: src/VX_sp_ram.sv:130:29
								ram[addr] <= wdata;
							if (read)
								// Trace: src/VX_sp_ram.sv:133:29
								rdata_r <= ram[addr];
						end
						// Trace: src/VX_sp_ram.sv:136:21
						assign rdata = rdata_r;
					end
				end
				else if (RDW_MODE == "N") begin : g_no_change
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:140:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:143:13
								initial begin
									// Trace: src/VX_sp_ram.sv:143:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:145:13
								initial begin
									// Trace: src/VX_sp_ram.sv:146:17
									begin : sv2v_autoblock_7
										// Trace: src/VX_sp_ram.sv:146:22
										integer i;
										// Trace: src/VX_sp_ram.sv:146:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:147:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:152:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:153:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:154:29
							if (write)
								// Trace: src/VX_sp_ram.sv:155:33
								begin : sv2v_autoblock_8
									// Trace: src/VX_sp_ram.sv:155:38
									integer i;
									// Trace: src/VX_sp_ram.sv:155:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:156:37
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:157:41
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							else if (read)
								// Trace: src/VX_sp_ram.sv:162:29
								rdata_r <= ram[addr];
						// Trace: src/VX_sp_ram.sv:165:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:167:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:170:13
								initial begin
									// Trace: src/VX_sp_ram.sv:170:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:172:13
								initial begin
									// Trace: src/VX_sp_ram.sv:173:17
									begin : sv2v_autoblock_9
										// Trace: src/VX_sp_ram.sv:173:22
										integer i;
										// Trace: src/VX_sp_ram.sv:173:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:174:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:179:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:180:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:181:25
							if (write)
								// Trace: src/VX_sp_ram.sv:182:29
								ram[addr] <= wdata;
							else if (read)
								// Trace: src/VX_sp_ram.sv:185:29
								rdata_r <= ram[addr];
						// Trace: src/VX_sp_ram.sv:188:21
						assign rdata = rdata_r;
					end
				end
			end
			else begin : g_auto
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:194:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:197:13
								initial begin
									// Trace: src/VX_sp_ram.sv:197:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:199:13
								initial begin
									// Trace: src/VX_sp_ram.sv:200:17
									begin : sv2v_autoblock_10
										// Trace: src/VX_sp_ram.sv:200:22
										integer i;
										// Trace: src/VX_sp_ram.sv:200:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:201:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:206:21
						reg [ADDRW - 1:0] addr_r;
						// Trace: src/VX_sp_ram.sv:207:21
						always @(posedge clk) begin
							// Trace: src/VX_sp_ram.sv:208:29
							if (write)
								// Trace: src/VX_sp_ram.sv:209:33
								begin : sv2v_autoblock_11
									// Trace: src/VX_sp_ram.sv:209:38
									integer i;
									// Trace: src/VX_sp_ram.sv:209:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:210:37
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:211:41
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							if (read)
								// Trace: src/VX_sp_ram.sv:216:29
								addr_r <= addr;
						end
						// Trace: src/VX_sp_ram.sv:219:21
						assign rdata = ram[addr_r];
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:221:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:224:13
								initial begin
									// Trace: src/VX_sp_ram.sv:224:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:226:13
								initial begin
									// Trace: src/VX_sp_ram.sv:227:17
									begin : sv2v_autoblock_12
										// Trace: src/VX_sp_ram.sv:227:22
										integer i;
										// Trace: src/VX_sp_ram.sv:227:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:228:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:233:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:234:21
						always @(posedge clk) begin
							// Trace: src/VX_sp_ram.sv:235:25
							if (write)
								// Trace: src/VX_sp_ram.sv:236:29
								ram[addr] <= wdata;
							if (read) begin
								begin
									// Trace: src/VX_sp_ram.sv:239:29
									if (write)
										// Trace: src/VX_sp_ram.sv:240:33
										rdata_r <= wdata;
									else
										// Trace: src/VX_sp_ram.sv:242:33
										rdata_r <= ram[addr];
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:246:21
						assign rdata = rdata_r;
					end
				end
				else if (RDW_MODE == "R") begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:250:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:253:13
								initial begin
									// Trace: src/VX_sp_ram.sv:253:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:255:13
								initial begin
									// Trace: src/VX_sp_ram.sv:256:17
									begin : sv2v_autoblock_13
										// Trace: src/VX_sp_ram.sv:256:22
										integer i;
										// Trace: src/VX_sp_ram.sv:256:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:257:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:262:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:263:21
						always @(posedge clk) begin
							// Trace: src/VX_sp_ram.sv:264:29
							if (write)
								// Trace: src/VX_sp_ram.sv:265:33
								begin : sv2v_autoblock_14
									// Trace: src/VX_sp_ram.sv:265:38
									integer i;
									// Trace: src/VX_sp_ram.sv:265:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:266:37
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:267:41
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							if (read)
								// Trace: src/VX_sp_ram.sv:272:29
								rdata_r <= ram[addr];
						end
						// Trace: src/VX_sp_ram.sv:275:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:277:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:280:13
								initial begin
									// Trace: src/VX_sp_ram.sv:280:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:282:13
								initial begin
									// Trace: src/VX_sp_ram.sv:283:17
									begin : sv2v_autoblock_15
										// Trace: src/VX_sp_ram.sv:283:22
										integer i;
										// Trace: src/VX_sp_ram.sv:283:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:284:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:289:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:290:21
						always @(posedge clk) begin
							// Trace: src/VX_sp_ram.sv:291:25
							if (write)
								// Trace: src/VX_sp_ram.sv:292:29
								ram[addr] <= wdata;
							if (read)
								// Trace: src/VX_sp_ram.sv:295:29
								rdata_r <= ram[addr];
						end
						// Trace: src/VX_sp_ram.sv:298:21
						assign rdata = rdata_r;
					end
				end
				else if (RDW_MODE == "N") begin : g_no_change
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:302:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:305:13
								initial begin
									// Trace: src/VX_sp_ram.sv:305:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:307:13
								initial begin
									// Trace: src/VX_sp_ram.sv:308:17
									begin : sv2v_autoblock_16
										// Trace: src/VX_sp_ram.sv:308:22
										integer i;
										// Trace: src/VX_sp_ram.sv:308:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:309:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:314:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:315:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:316:29
							if (write)
								// Trace: src/VX_sp_ram.sv:317:33
								begin : sv2v_autoblock_17
									// Trace: src/VX_sp_ram.sv:317:38
									integer i;
									// Trace: src/VX_sp_ram.sv:317:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:318:37
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:319:41
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							else if (read)
								// Trace: src/VX_sp_ram.sv:324:29
								rdata_r <= ram[addr];
						// Trace: src/VX_sp_ram.sv:327:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:329:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:332:13
								initial begin
									// Trace: src/VX_sp_ram.sv:332:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:334:13
								initial begin
									// Trace: src/VX_sp_ram.sv:335:17
									begin : sv2v_autoblock_18
										// Trace: src/VX_sp_ram.sv:335:22
										integer i;
										// Trace: src/VX_sp_ram.sv:335:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:336:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:341:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_sp_ram.sv:342:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:343:25
							if (write)
								// Trace: src/VX_sp_ram.sv:344:29
								ram[addr] <= wdata;
							else if (read)
								// Trace: src/VX_sp_ram.sv:347:29
								rdata_r <= ram[addr];
						// Trace: src/VX_sp_ram.sv:350:21
						assign rdata = rdata_r;
					end
				end
			end
		end
		else begin : g_async
			if (FORCE_BRAM) begin : g_bram
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:358:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:361:13
								initial begin
									// Trace: src/VX_sp_ram.sv:361:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:363:13
								initial begin
									// Trace: src/VX_sp_ram.sv:364:17
									begin : sv2v_autoblock_19
										// Trace: src/VX_sp_ram.sv:364:22
										integer i;
										// Trace: src/VX_sp_ram.sv:364:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:365:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:370:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:371:29
							if (write)
								// Trace: src/VX_sp_ram.sv:372:33
								begin : sv2v_autoblock_20
									// Trace: src/VX_sp_ram.sv:372:38
									integer i;
									// Trace: src/VX_sp_ram.sv:372:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:373:37
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:374:41
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_sp_ram.sv:379:21
						assign rdata = ram[addr];
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:381:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:384:13
								initial begin
									// Trace: src/VX_sp_ram.sv:384:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:386:13
								initial begin
									// Trace: src/VX_sp_ram.sv:387:17
									begin : sv2v_autoblock_21
										// Trace: src/VX_sp_ram.sv:387:22
										integer i;
										// Trace: src/VX_sp_ram.sv:387:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:388:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:393:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:394:25
							if (write)
								// Trace: src/VX_sp_ram.sv:395:29
								ram[addr] <= wdata;
						// Trace: src/VX_sp_ram.sv:398:21
						assign rdata = ram[addr];
					end
				end
				else begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:402:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:405:13
								initial begin
									// Trace: src/VX_sp_ram.sv:405:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:407:13
								initial begin
									// Trace: src/VX_sp_ram.sv:408:17
									begin : sv2v_autoblock_22
										// Trace: src/VX_sp_ram.sv:408:22
										integer i;
										// Trace: src/VX_sp_ram.sv:408:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:409:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:414:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:415:29
							if (write)
								// Trace: src/VX_sp_ram.sv:416:33
								begin : sv2v_autoblock_23
									// Trace: src/VX_sp_ram.sv:416:38
									integer i;
									// Trace: src/VX_sp_ram.sv:416:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:417:37
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:418:41
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_sp_ram.sv:423:21
						assign rdata = ram[addr];
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:425:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:428:13
								initial begin
									// Trace: src/VX_sp_ram.sv:428:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:430:13
								initial begin
									// Trace: src/VX_sp_ram.sv:431:17
									begin : sv2v_autoblock_24
										// Trace: src/VX_sp_ram.sv:431:22
										integer i;
										// Trace: src/VX_sp_ram.sv:431:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:432:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:437:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:438:25
							if (write)
								// Trace: src/VX_sp_ram.sv:439:29
								ram[addr] <= wdata;
						// Trace: src/VX_sp_ram.sv:442:21
						assign rdata = ram[addr];
					end
				end
			end
			else begin : g_auto
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:448:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:451:13
								initial begin
									// Trace: src/VX_sp_ram.sv:451:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:453:13
								initial begin
									// Trace: src/VX_sp_ram.sv:454:17
									begin : sv2v_autoblock_25
										// Trace: src/VX_sp_ram.sv:454:22
										integer i;
										// Trace: src/VX_sp_ram.sv:454:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:455:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:460:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:461:29
							if (write)
								// Trace: src/VX_sp_ram.sv:462:33
								begin : sv2v_autoblock_26
									// Trace: src/VX_sp_ram.sv:462:38
									integer i;
									// Trace: src/VX_sp_ram.sv:462:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:463:37
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:464:41
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_sp_ram.sv:469:21
						assign rdata = ram[addr];
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:471:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:474:13
								initial begin
									// Trace: src/VX_sp_ram.sv:474:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:476:13
								initial begin
									// Trace: src/VX_sp_ram.sv:477:17
									begin : sv2v_autoblock_27
										// Trace: src/VX_sp_ram.sv:477:22
										integer i;
										// Trace: src/VX_sp_ram.sv:477:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:478:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:483:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:484:25
							if (write)
								// Trace: src/VX_sp_ram.sv:485:29
								ram[addr] <= wdata;
						// Trace: src/VX_sp_ram.sv:488:21
						assign rdata = ram[addr];
					end
				end
				else begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_sp_ram.sv:492:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:495:13
								initial begin
									// Trace: src/VX_sp_ram.sv:495:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:497:13
								initial begin
									// Trace: src/VX_sp_ram.sv:498:17
									begin : sv2v_autoblock_28
										// Trace: src/VX_sp_ram.sv:498:22
										integer i;
										// Trace: src/VX_sp_ram.sv:498:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:499:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:504:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:505:29
							if (write)
								// Trace: src/VX_sp_ram.sv:506:33
								begin : sv2v_autoblock_29
									// Trace: src/VX_sp_ram.sv:506:38
									integer i;
									// Trace: src/VX_sp_ram.sv:506:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_sp_ram.sv:507:37
											if (wren[i])
												// Trace: src/VX_sp_ram.sv:508:41
												ram[addr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_sp_ram.sv:513:21
						assign rdata = ram[addr];
					end
					else begin : g_no_wren
						// Trace: src/VX_sp_ram.sv:515:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_sp_ram.sv:518:13
								initial begin
									// Trace: src/VX_sp_ram.sv:518:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_sp_ram.sv:520:13
								initial begin
									// Trace: src/VX_sp_ram.sv:521:17
									begin : sv2v_autoblock_30
										// Trace: src/VX_sp_ram.sv:521:22
										integer i;
										// Trace: src/VX_sp_ram.sv:521:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_sp_ram.sv:522:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_sp_ram.sv:527:21
						always @(posedge clk)
							// Trace: src/VX_sp_ram.sv:528:25
							if (write)
								// Trace: src/VX_sp_ram.sv:529:29
								ram[addr] <= wdata;
						// Trace: src/VX_sp_ram.sv:532:21
						assign rdata = ram[addr];
					end
				end
			end
		end
	endgenerate
endmodule
module VX_transpose (
	data_in,
	data_out
);
	// Trace: src/VX_transpose.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_transpose.sv:3:15
	parameter N = 1;
	// Trace: src/VX_transpose.sv:4:15
	parameter M = 1;
	// Trace: src/VX_transpose.sv:6:5
	input wire [((N * M) * DATAW) - 1:0] data_in;
	// Trace: src/VX_transpose.sv:7:5
	output wire [((M * N) * DATAW) - 1:0] data_out;
	// Trace: src/VX_transpose.sv:9:5
	genvar _gv_i_126;
	generate
		for (_gv_i_126 = 0; _gv_i_126 < N; _gv_i_126 = _gv_i_126 + 1) begin : g_i
			localparam i = _gv_i_126;
			genvar _gv_j_14;
			for (_gv_j_14 = 0; _gv_j_14 < M; _gv_j_14 = _gv_j_14 + 1) begin : g_j
				localparam j = _gv_j_14;
				// Trace: src/VX_transpose.sv:11:13
				assign data_out[((j * N) + i) * DATAW+:DATAW] = data_in[((i * M) + j) * DATAW+:DATAW];
			end
		end
	endgenerate
endmodule
// removed module with interface ports: VX_decode
// removed module with interface ports: VX_mem_unit
// removed interface: VX_commit_csr_if
module VX_demux (
	sel_in,
	data_in,
	data_out
);
	// Trace: src/VX_demux.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_demux.sv:3:15
	parameter N = 0;
	// Trace: src/VX_demux.sv:4:15
	parameter MODEL = 0;
	// Trace: src/VX_demux.sv:5:15
	parameter LN = (N > 1 ? $clog2(N) : 1);
	// Trace: src/VX_demux.sv:7:5
	input wire [LN - 1:0] sel_in;
	// Trace: src/VX_demux.sv:8:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_demux.sv:9:5
	output wire [(N * DATAW) - 1:0] data_out;
	// Trace: src/VX_demux.sv:11:5
	function automatic [(N * DATAW) - 1:0] sv2v_cast_3AE7C;
		input reg [(N * DATAW) - 1:0] inp;
		sv2v_cast_3AE7C = inp;
	endfunction
	generate
		if (N > 1) begin : g_demux
			// Trace: src/VX_demux.sv:12:9
			reg [(N * DATAW) - 1:0] shift;
			if (MODEL == 1) begin : g_model1
				// Trace: src/VX_demux.sv:14:13
				always @(*) begin
					// Trace: src/VX_demux.sv:15:17
					shift = 1'sb0;
					// Trace: src/VX_demux.sv:16:17
					shift[sel_in * DATAW+:DATAW] = {DATAW {1'b1}};
				end
			end
			else begin : g_model0
				// Trace: src/VX_demux.sv:19:13
				wire [N * DATAW:1] sv2v_tmp_6BA10;
				assign sv2v_tmp_6BA10 = sv2v_cast_3AE7C({DATAW {1'b1}}) << (sel_in * DATAW);
				always @(*) shift = sv2v_tmp_6BA10;
			end
			// Trace: src/VX_demux.sv:21:9
			assign data_out = {N {data_in}} & shift;
		end
		else begin : g_passthru
			// Trace: src/VX_demux.sv:23:9
			assign data_out = data_in;
		end
	endgenerate
endmodule
module VX_rr_arbiter (
	clk,
	reset,
	requests,
	grant_index,
	grant_onehot,
	grant_valid,
	grant_ready
);
	// Trace: src/VX_rr_arbiter.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_rr_arbiter.sv:3:15
	parameter MODEL = 1;
	// Trace: src/VX_rr_arbiter.sv:4:15
	parameter LOG_NUM_REQS = (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1);
	// Trace: src/VX_rr_arbiter.sv:5:15
	parameter STICKY = 0;
	// Trace: src/VX_rr_arbiter.sv:6:15
	parameter LUT_OPT = 0;
	// Trace: src/VX_rr_arbiter.sv:8:5
	input wire clk;
	// Trace: src/VX_rr_arbiter.sv:9:5
	input wire reset;
	// Trace: src/VX_rr_arbiter.sv:10:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: src/VX_rr_arbiter.sv:11:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: src/VX_rr_arbiter.sv:12:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: src/VX_rr_arbiter.sv:13:5
	output wire grant_valid;
	// Trace: src/VX_rr_arbiter.sv:14:5
	input wire grant_ready;
	// Trace: src/VX_rr_arbiter.sv:16:5
	function automatic signed [LOG_NUM_REQS - 1:0] sv2v_cast_76B5F_signed;
		input reg signed [LOG_NUM_REQS - 1:0] inp;
		sv2v_cast_76B5F_signed = inp;
	endfunction
	generate
		if (NUM_REQS == 1) begin : g_passthru
			// Trace: src/VX_rr_arbiter.sv:17:9
			assign grant_index = 1'sb0;
			// Trace: src/VX_rr_arbiter.sv:18:9
			assign grant_onehot = requests;
			// Trace: src/VX_rr_arbiter.sv:19:9
			assign grant_valid = requests[0];
		end
		else if (LUT_OPT && (NUM_REQS == 2)) begin : g_lut2
			// Trace: src/VX_rr_arbiter.sv:21:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:22:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:23:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:24:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:25:13
				casez ({state, requests})
					3'b001, 3'b1z1: begin
						// Trace: src/VX_rr_arbiter.sv:27:28
						grant_onehot_w = 2'b01;
						// Trace: src/VX_rr_arbiter.sv:27:52
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					3'b01z, 3'b110: begin
						// Trace: src/VX_rr_arbiter.sv:29:28
						grant_onehot_w = 2'b10;
						// Trace: src/VX_rr_arbiter.sv:29:52
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:30:28
						grant_onehot_w = 2'b00;
						// Trace: src/VX_rr_arbiter.sv:30:52
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:33:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:34:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:35:17
					state <= 1'sb0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_rr_arbiter.sv:37:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:40:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:41:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:42:9
			assign grant_valid = |requests;
		end
		else if (LUT_OPT && (NUM_REQS == 3)) begin : g_lut3
			// Trace: src/VX_rr_arbiter.sv:44:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:45:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:46:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:47:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:48:13
				casez ({state, requests})
					5'b00001, 5'b010z1, 5'b10zz1: begin
						// Trace: src/VX_rr_arbiter.sv:51:30
						grant_onehot_w = 3'b001;
						// Trace: src/VX_rr_arbiter.sv:51:55
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					5'b00z1z, 5'b01010, 5'b10z10: begin
						// Trace: src/VX_rr_arbiter.sv:54:30
						grant_onehot_w = 3'b010;
						// Trace: src/VX_rr_arbiter.sv:54:55
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					5'b0010z, 5'b011zz, 5'b10100: begin
						// Trace: src/VX_rr_arbiter.sv:57:30
						grant_onehot_w = 3'b100;
						// Trace: src/VX_rr_arbiter.sv:57:55
						grant_index_w = sv2v_cast_76B5F_signed(2);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:58:30
						grant_onehot_w = 3'b000;
						// Trace: src/VX_rr_arbiter.sv:58:55
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:61:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:62:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:63:17
					state <= 1'sb0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_rr_arbiter.sv:65:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:68:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:69:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:70:9
			assign grant_valid = |requests;
		end
		else if (LUT_OPT && (NUM_REQS == 4)) begin : g_lut4
			// Trace: src/VX_rr_arbiter.sv:72:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:73:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:74:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:75:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:76:13
				casez ({state, requests})
					6'b000001, 6'b0100z1, 6'b100zz1, 6'b11zzz1: begin
						// Trace: src/VX_rr_arbiter.sv:80:31
						grant_onehot_w = 4'b0001;
						// Trace: src/VX_rr_arbiter.sv:80:57
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					6'b00zz1z, 6'b010010, 6'b100z10, 6'b11zz10: begin
						// Trace: src/VX_rr_arbiter.sv:84:31
						grant_onehot_w = 4'b0010;
						// Trace: src/VX_rr_arbiter.sv:84:57
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					6'b00z10z, 6'b01z1zz, 6'b100100, 6'b11z100: begin
						// Trace: src/VX_rr_arbiter.sv:88:31
						grant_onehot_w = 4'b0100;
						// Trace: src/VX_rr_arbiter.sv:88:57
						grant_index_w = sv2v_cast_76B5F_signed(2);
					end
					6'b00100z, 6'b0110zz, 6'b101zzz, 6'b111000: begin
						// Trace: src/VX_rr_arbiter.sv:92:31
						grant_onehot_w = 4'b1000;
						// Trace: src/VX_rr_arbiter.sv:92:57
						grant_index_w = sv2v_cast_76B5F_signed(3);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:93:31
						grant_onehot_w = 4'b0000;
						// Trace: src/VX_rr_arbiter.sv:93:57
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:96:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:97:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:98:17
					state <= 1'sb0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_rr_arbiter.sv:100:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:103:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:104:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:105:9
			assign grant_valid = |requests;
		end
		else if (LUT_OPT && (NUM_REQS == 5)) begin : g_lut5
			// Trace: src/VX_rr_arbiter.sv:107:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:108:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:109:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:110:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:111:13
				casez ({state, requests})
					8'b00000001, 8'b001000z1, 8'b01000zz1, 8'b0110zzz1, 8'b100zzzz1: begin
						// Trace: src/VX_rr_arbiter.sv:116:33
						grant_onehot_w = 5'b00001;
						// Trace: src/VX_rr_arbiter.sv:116:60
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					8'b000zzz1z, 8'b00100010, 8'b01000z10, 8'b0110zz10, 8'b100zzz10: begin
						// Trace: src/VX_rr_arbiter.sv:121:33
						grant_onehot_w = 5'b00010;
						// Trace: src/VX_rr_arbiter.sv:121:60
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					8'b000zz10z, 8'b001zz1zz, 8'b01000100, 8'b0110z100, 8'b100zz100: begin
						// Trace: src/VX_rr_arbiter.sv:126:33
						grant_onehot_w = 5'b00100;
						// Trace: src/VX_rr_arbiter.sv:126:60
						grant_index_w = sv2v_cast_76B5F_signed(2);
					end
					8'b000z100z, 8'b001z10zz, 8'b010z1zzz, 8'b01101000, 8'b100z1000: begin
						// Trace: src/VX_rr_arbiter.sv:131:33
						grant_onehot_w = 5'b01000;
						// Trace: src/VX_rr_arbiter.sv:131:60
						grant_index_w = sv2v_cast_76B5F_signed(3);
					end
					8'b0001000z, 8'b001100zz, 8'b01010zzz, 8'b0111zzzz, 8'b10010000: begin
						// Trace: src/VX_rr_arbiter.sv:136:33
						grant_onehot_w = 5'b10000;
						// Trace: src/VX_rr_arbiter.sv:136:60
						grant_index_w = sv2v_cast_76B5F_signed(4);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:137:33
						grant_onehot_w = 5'b00000;
						// Trace: src/VX_rr_arbiter.sv:137:60
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:140:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:141:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:142:17
					state <= 1'sb0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_rr_arbiter.sv:144:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:147:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:148:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:149:9
			assign grant_valid = |requests;
		end
		else if (LUT_OPT && (NUM_REQS == 6)) begin : g_lut6
			// Trace: src/VX_rr_arbiter.sv:151:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:152:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:153:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:154:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:155:13
				casez ({state, requests})
					9'b000000001, 9'b0010000z1, 9'b010000zz1, 9'b01100zzz1, 9'b1000zzzz1, 9'b101zzzzz1: begin
						// Trace: src/VX_rr_arbiter.sv:161:34
						grant_onehot_w = 6'b000001;
						// Trace: src/VX_rr_arbiter.sv:161:62
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					9'b000zzzz1z, 9'b001000010, 9'b010000z10, 9'b01100zz10, 9'b1000zzz10, 9'b101zzzz10: begin
						// Trace: src/VX_rr_arbiter.sv:167:34
						grant_onehot_w = 6'b000010;
						// Trace: src/VX_rr_arbiter.sv:167:62
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					9'b000zzz10z, 9'b001zzz1zz, 9'b010000100, 9'b01100z100, 9'b1000zz100, 9'b101zzz100: begin
						// Trace: src/VX_rr_arbiter.sv:173:34
						grant_onehot_w = 6'b000100;
						// Trace: src/VX_rr_arbiter.sv:173:62
						grant_index_w = sv2v_cast_76B5F_signed(2);
					end
					9'b000zz100z, 9'b001zz10zz, 9'b010zz1zzz, 9'b011001000, 9'b1000z1000, 9'b101zz1000: begin
						// Trace: src/VX_rr_arbiter.sv:179:34
						grant_onehot_w = 6'b001000;
						// Trace: src/VX_rr_arbiter.sv:179:62
						grant_index_w = sv2v_cast_76B5F_signed(3);
					end
					9'b000z1000z, 9'b001z100zz, 9'b010z10zzz, 9'b011z1zzzz, 9'b100010000, 9'b101z10000: begin
						// Trace: src/VX_rr_arbiter.sv:185:34
						grant_onehot_w = 6'b010000;
						// Trace: src/VX_rr_arbiter.sv:185:62
						grant_index_w = sv2v_cast_76B5F_signed(4);
					end
					9'b00010000z, 9'b0011000zz, 9'b010100zzz, 9'b01110zzzz, 9'b1001zzzzz, 9'b101100000: begin
						// Trace: src/VX_rr_arbiter.sv:191:34
						grant_onehot_w = 6'b100000;
						// Trace: src/VX_rr_arbiter.sv:191:62
						grant_index_w = sv2v_cast_76B5F_signed(5);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:192:34
						grant_onehot_w = 6'b000000;
						// Trace: src/VX_rr_arbiter.sv:192:62
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:195:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:196:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:197:17
					state <= 1'sb0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_rr_arbiter.sv:199:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:202:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:203:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:204:9
			assign grant_valid = |requests;
		end
		else if (LUT_OPT && (NUM_REQS == 7)) begin : g_lut7
			// Trace: src/VX_rr_arbiter.sv:206:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:207:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:208:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:209:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:210:13
				casez ({state, requests})
					10'b0000000001, 10'b00100000z1, 10'b0100000zz1, 10'b011000zzz1, 10'b100000zzz1, 10'b10100zzzz1, 10'b110zzzzzz1: begin
						// Trace: src/VX_rr_arbiter.sv:217:36
						grant_onehot_w = 7'b0000001;
						// Trace: src/VX_rr_arbiter.sv:217:65
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					10'b000zzzzz1z, 10'b0010000010, 10'b0100000z10, 10'b011000zz10, 10'b10000zzz10, 10'b1010zzzz10, 10'b110zzzzz10: begin
						// Trace: src/VX_rr_arbiter.sv:224:36
						grant_onehot_w = 7'b0000010;
						// Trace: src/VX_rr_arbiter.sv:224:65
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					10'b000zzzz10z, 10'b001zzzz1zz, 10'b0100000100, 10'b011000z100, 10'b10000zz100, 10'b1010zzz100, 10'b110zzzz100: begin
						// Trace: src/VX_rr_arbiter.sv:231:36
						grant_onehot_w = 7'b0000100;
						// Trace: src/VX_rr_arbiter.sv:231:65
						grant_index_w = sv2v_cast_76B5F_signed(2);
					end
					10'b000zzz100z, 10'b001zzz10zz, 10'b010zzz1zzz, 10'b0110001000, 10'b10000z1000, 10'b1010zz1000, 10'b110zzz1000: begin
						// Trace: src/VX_rr_arbiter.sv:238:36
						grant_onehot_w = 7'b0001000;
						// Trace: src/VX_rr_arbiter.sv:238:65
						grant_index_w = sv2v_cast_76B5F_signed(3);
					end
					10'b000zz1000z, 10'b001zz100zz, 10'b010zz10zzz, 10'b011zz1zzzz, 10'b1000010000, 10'b1010z10000, 10'b110zz10000: begin
						// Trace: src/VX_rr_arbiter.sv:245:36
						grant_onehot_w = 7'b0010000;
						// Trace: src/VX_rr_arbiter.sv:245:65
						grant_index_w = sv2v_cast_76B5F_signed(4);
					end
					10'b000z10000z, 10'b001z1000zz, 10'b010z100zzz, 10'b011z10zzzz, 10'b100z1zzzzz, 10'b1010100000, 10'b110z100000: begin
						// Trace: src/VX_rr_arbiter.sv:252:36
						grant_onehot_w = 7'b0100000;
						// Trace: src/VX_rr_arbiter.sv:252:65
						grant_index_w = sv2v_cast_76B5F_signed(5);
					end
					10'b000100000z, 10'b00110000zz, 10'b0101000zzz, 10'b011100zzzz, 10'b10010zzzzz, 10'b1011zzzzzz, 10'b1101000000: begin
						// Trace: src/VX_rr_arbiter.sv:259:36
						grant_onehot_w = 7'b1000000;
						// Trace: src/VX_rr_arbiter.sv:259:65
						grant_index_w = sv2v_cast_76B5F_signed(6);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:260:35
						grant_onehot_w = 7'b0000000;
						// Trace: src/VX_rr_arbiter.sv:260:64
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:263:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:264:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:265:17
					state <= 1'sb0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_rr_arbiter.sv:267:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:270:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:271:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:272:9
			assign grant_valid = |requests;
		end
		else if (LUT_OPT && (NUM_REQS == 8)) begin : g_lut8
			// Trace: src/VX_rr_arbiter.sv:274:9
			reg [LOG_NUM_REQS - 1:0] grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:275:9
			reg [NUM_REQS - 1:0] grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:276:9
			reg [LOG_NUM_REQS - 1:0] state;
			// Trace: src/VX_rr_arbiter.sv:277:9
			always @(*)
				// Trace: src/VX_rr_arbiter.sv:278:13
				casez ({state, requests})
					11'b00000000001, 11'b001000000z1, 11'b01000000zz1, 11'b0110000zzz1, 11'b100000zzzz1, 11'b10100zzzzz1, 11'b1100zzzzzz1, 11'b111zzzzzzz1: begin
						// Trace: src/VX_rr_arbiter.sv:286:37
						grant_onehot_w = 8'b00000001;
						// Trace: src/VX_rr_arbiter.sv:286:67
						grant_index_w = sv2v_cast_76B5F_signed(0);
					end
					11'b000zzzzzz1z, 11'b00100000010, 11'b01000000z10, 11'b0110000zz10, 11'b100000zzz10, 11'b10100zzzz10, 11'b1100zzzzz10, 11'b111zzzzzz10: begin
						// Trace: src/VX_rr_arbiter.sv:294:37
						grant_onehot_w = 8'b00000010;
						// Trace: src/VX_rr_arbiter.sv:294:67
						grant_index_w = sv2v_cast_76B5F_signed(1);
					end
					11'b000zzzzz10z, 11'b001zzzzz1zz, 11'b01000000100, 11'b0110000z100, 11'b100000zz100, 11'b10100zzz100, 11'b1100zzzz100, 11'b111zzzzz100: begin
						// Trace: src/VX_rr_arbiter.sv:302:37
						grant_onehot_w = 8'b00000100;
						// Trace: src/VX_rr_arbiter.sv:302:67
						grant_index_w = sv2v_cast_76B5F_signed(2);
					end
					11'b000zzzz100z, 11'b001zzzz10zz, 11'b010zzzz1zzz, 11'b01100001000, 11'b100000z1000, 11'b10100zz1000, 11'b1100zzz1000, 11'b111zzzz1000: begin
						// Trace: src/VX_rr_arbiter.sv:310:37
						grant_onehot_w = 8'b00001000;
						// Trace: src/VX_rr_arbiter.sv:310:67
						grant_index_w = sv2v_cast_76B5F_signed(3);
					end
					11'b000zzz1000z, 11'b001zzz100zz, 11'b010zzz10zzz, 11'b011zzz1zzzz, 11'b10000010000, 11'b10100z10000, 11'b1100zz10000, 11'b111zzz10000: begin
						// Trace: src/VX_rr_arbiter.sv:318:37
						grant_onehot_w = 8'b00010000;
						// Trace: src/VX_rr_arbiter.sv:318:67
						grant_index_w = sv2v_cast_76B5F_signed(4);
					end
					11'b000zz10000z, 11'b001zz1000zz, 11'b010zz100zzz, 11'b011zz10zzzz, 11'b100zz1zzzzz, 11'b10100100000, 11'b1100z100000, 11'b111zz100000: begin
						// Trace: src/VX_rr_arbiter.sv:326:37
						grant_onehot_w = 8'b00100000;
						// Trace: src/VX_rr_arbiter.sv:326:67
						grant_index_w = sv2v_cast_76B5F_signed(5);
					end
					11'b000z100000z, 11'b001z10000zz, 11'b010z1000zzz, 11'b011z100zzzz, 11'b100z10zzzzz, 11'b101z1zzzzzz, 11'b11001000000, 11'b111z1000000: begin
						// Trace: src/VX_rr_arbiter.sv:334:37
						grant_onehot_w = 8'b01000000;
						// Trace: src/VX_rr_arbiter.sv:334:67
						grant_index_w = sv2v_cast_76B5F_signed(6);
					end
					11'b0001000000z, 11'b001100000zz, 11'b01010000zzz, 11'b0111000zzzz, 11'b100100zzzzz, 11'b10110zzzzzz, 11'b1101zzzzzzz, 11'b11110000000: begin
						// Trace: src/VX_rr_arbiter.sv:342:37
						grant_onehot_w = 8'b10000000;
						// Trace: src/VX_rr_arbiter.sv:342:67
						grant_index_w = sv2v_cast_76B5F_signed(7);
					end
					default: begin
						// Trace: src/VX_rr_arbiter.sv:343:37
						grant_onehot_w = 8'b00000000;
						// Trace: src/VX_rr_arbiter.sv:343:67
						grant_index_w = 1'sbx;
					end
				endcase
			// Trace: src/VX_rr_arbiter.sv:346:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:347:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:348:17
					state <= 1'sb0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_rr_arbiter.sv:350:17
					state <= grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:353:9
			assign grant_index = grant_index_w;
			// Trace: src/VX_rr_arbiter.sv:354:9
			assign grant_onehot = grant_onehot_w;
			// Trace: src/VX_rr_arbiter.sv:355:9
			assign grant_valid = |requests;
		end
		else if (MODEL == 1) begin : g_model1
			// Trace: src/VX_rr_arbiter.sv:357:9
			wire [NUM_REQS - 1:0] masked_pri_reqs;
			wire [NUM_REQS - 1:0] unmasked_pri_reqs;
			// Trace: src/VX_rr_arbiter.sv:358:9
			reg [NUM_REQS - 1:0] reqs_mask;
			// Trace: src/VX_rr_arbiter.sv:359:9
			wire [NUM_REQS - 1:0] masked_reqs = requests & reqs_mask;
			// Trace: src/VX_rr_arbiter.sv:360:9
			assign masked_pri_reqs[0] = 1'b0;
			genvar _gv_i_131;
			for (_gv_i_131 = 1; _gv_i_131 < NUM_REQS; _gv_i_131 = _gv_i_131 + 1) begin : g_masked_pri_reqs
				localparam i = _gv_i_131;
				// Trace: src/VX_rr_arbiter.sv:362:13
				assign masked_pri_reqs[i] = masked_pri_reqs[i - 1] | masked_reqs[i - 1];
			end
			// Trace: src/VX_rr_arbiter.sv:364:9
			assign unmasked_pri_reqs[0] = 1'b0;
			genvar _gv_i_132;
			for (_gv_i_132 = 1; _gv_i_132 < NUM_REQS; _gv_i_132 = _gv_i_132 + 1) begin : g_unmasked_pri_reqs
				localparam i = _gv_i_132;
				// Trace: src/VX_rr_arbiter.sv:366:13
				assign unmasked_pri_reqs[i] = unmasked_pri_reqs[i - 1] | requests[i - 1];
			end
			// Trace: src/VX_rr_arbiter.sv:368:9
			wire [NUM_REQS - 1:0] grant_masked = masked_reqs & ~masked_pri_reqs;
			// Trace: src/VX_rr_arbiter.sv:369:9
			wire [NUM_REQS - 1:0] grant_unmasked = requests & ~unmasked_pri_reqs;
			// Trace: src/VX_rr_arbiter.sv:370:9
			wire has_masked_reqs = |masked_reqs;
			// Trace: src/VX_rr_arbiter.sv:371:9
			wire has_unmasked_reqs = |requests;
			// Trace: src/VX_rr_arbiter.sv:372:9
			reg [NUM_REQS - 1:0] prev_grant;
			// Trace: src/VX_rr_arbiter.sv:373:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:374:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:375:17
					prev_grant <= 1'sb0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_rr_arbiter.sv:377:17
					prev_grant <= grant_onehot;
			// Trace: src/VX_rr_arbiter.sv:380:9
			wire retain_grant = (STICKY != 0) && |(prev_grant & requests);
			// Trace: src/VX_rr_arbiter.sv:381:9
			wire [NUM_REQS - 1:0] grant = (has_masked_reqs ? grant_masked : grant_unmasked);
			// Trace: src/VX_rr_arbiter.sv:382:9
			wire [NUM_REQS - 1:0] grant_w = (retain_grant ? prev_grant : grant);
			// Trace: src/VX_rr_arbiter.sv:383:9
			assign grant_onehot = grant_w;
			// Trace: src/VX_rr_arbiter.sv:384:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:385:7
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:386:5
					reqs_mask <= {NUM_REQS {1'b1}};
				else if ((grant_valid && grant_ready) && ~retain_grant) begin
					begin
						// Trace: src/VX_rr_arbiter.sv:388:5
						if (has_masked_reqs)
							// Trace: src/VX_rr_arbiter.sv:389:21
							reqs_mask <= masked_pri_reqs;
						else if (has_unmasked_reqs)
							// Trace: src/VX_rr_arbiter.sv:391:21
							reqs_mask <= unmasked_pri_reqs;
					end
				end
			// Trace: src/VX_rr_arbiter.sv:395:9
			wire grant_valid_w;
			// Trace: src/VX_rr_arbiter.sv:396:9
			VX_onehot_encoder #(.N(NUM_REQS)) onehot_encoder(
				.data_in(grant_w),
				.data_out(grant_index),
				.valid_out(grant_valid_w)
			);
			// Trace: src/VX_rr_arbiter.sv:403:9
			assign grant_valid = (STICKY != 0 ? |requests : grant_valid_w);
		end
		else if (MODEL == 2) begin : g_model2
			// Trace: src/VX_rr_arbiter.sv:405:9
			reg [(NUM_REQS * LOG_NUM_REQS) - 1:0] grant_table;
			// Trace: src/VX_rr_arbiter.sv:406:9
			reg [LOG_NUM_REQS - 1:0] state;
			genvar _gv_i_133;
			for (_gv_i_133 = 0; _gv_i_133 < NUM_REQS; _gv_i_133 = _gv_i_133 + 1) begin : g_grant_table
				localparam i = _gv_i_133;
				// Trace: src/VX_rr_arbiter.sv:408:13
				always @(*) begin
					// Trace: src/VX_rr_arbiter.sv:409:17
					grant_table[i * LOG_NUM_REQS+:LOG_NUM_REQS] = 1'sbx;
					// Trace: src/VX_rr_arbiter.sv:410:17
					begin : sv2v_autoblock_1
						// Trace: src/VX_rr_arbiter.sv:410:22
						integer j;
						// Trace: src/VX_rr_arbiter.sv:410:22
						for (j = NUM_REQS - 1; j >= 0; j = j - 1)
							begin
								// Trace: src/VX_rr_arbiter.sv:411:21
								if (requests[((i + j) + 1) % NUM_REQS])
									// Trace: src/VX_rr_arbiter.sv:412:25
									grant_table[i * LOG_NUM_REQS+:LOG_NUM_REQS] = sv2v_cast_76B5F_signed(((i + j) + 1) % NUM_REQS);
							end
					end
				end
			end
			// Trace: src/VX_rr_arbiter.sv:417:9
			always @(posedge clk)
				// Trace: src/VX_rr_arbiter.sv:418:13
				if (reset)
					// Trace: src/VX_rr_arbiter.sv:419:17
					state <= 0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_rr_arbiter.sv:421:17
					state <= grant_index;
			// Trace: src/VX_rr_arbiter.sv:424:9
			VX_demux #(
				.DATAW(1),
				.N(NUM_REQS)
			) grant_decoder(
				.sel_in(grant_index),
				.data_in(grant_valid),
				.data_out(grant_onehot)
			);
			// Trace: src/VX_rr_arbiter.sv:432:9
			assign grant_index = grant_table[state * LOG_NUM_REQS+:LOG_NUM_REQS];
			// Trace: src/VX_rr_arbiter.sv:433:9
			assign grant_valid = |requests;
		end
	endgenerate
endmodule
module VX_split_join (
	clk,
	reset,
	valid,
	wid,
	split,
	sjoin,
	stack_wid,
	join_valid,
	join_is_dvg,
	join_is_else,
	join_wid,
	join_tmask,
	join_pc,
	stack_ptr
);
	// removed import VX_gpu_pkg::*;
	// Trace: src/VX_split_join.sv:2:15
	parameter INSTANCE_ID = "";
	// Trace: src/VX_split_join.sv:3:15
	parameter OUT_REG = 0;
	// Trace: src/VX_split_join.sv:5:5
	input wire clk;
	// Trace: src/VX_split_join.sv:6:5
	input wire reset;
	// Trace: src/VX_split_join.sv:7:5
	input wire valid;
	// Trace: src/VX_split_join.sv:8:5
	localparam VX_gpu_pkg_NW_BITS = 2;
	localparam VX_gpu_pkg_NW_WIDTH = VX_gpu_pkg_NW_BITS;
	input wire [1:0] wid;
	// Trace: src/VX_split_join.sv:9:5
	localparam VX_gpu_pkg_PC_BITS = 30;
	// removed localparam type VX_gpu_pkg_split_t
	input wire [39:0] split;
	// Trace: src/VX_split_join.sv:10:5
	localparam VX_gpu_pkg_DV_STACK_SIZE = 3;
	localparam VX_gpu_pkg_DV_STACK_SIZEW = 2;
	// removed localparam type VX_gpu_pkg_join_t
	input wire [2:0] sjoin;
	// Trace: src/VX_split_join.sv:11:5
	input wire [1:0] stack_wid;
	// Trace: src/VX_split_join.sv:12:5
	output wire join_valid;
	// Trace: src/VX_split_join.sv:13:5
	output wire join_is_dvg;
	// Trace: src/VX_split_join.sv:14:5
	output wire join_is_else;
	// Trace: src/VX_split_join.sv:15:5
	output wire [1:0] join_wid;
	// Trace: src/VX_split_join.sv:16:5
	output wire [3:0] join_tmask;
	// Trace: src/VX_split_join.sv:17:5
	output wire [29:0] join_pc;
	// Trace: src/VX_split_join.sv:18:5
	output wire [1:0] stack_ptr;
	// Trace: src/VX_split_join.sv:20:5
	wire split_valid = valid && split[39];
	// Trace: src/VX_split_join.sv:21:5
	wire sjoin_valid = valid && sjoin[2];
	// Trace: src/VX_split_join.sv:22:5
	localparam VX_gpu_pkg_NT_BITS = 2;
	generate
		if (1) begin : g_enable
			// Trace: src/VX_split_join.sv:23:9
			wire [7:0] ipdom_wr_ptr;
			// Trace: src/VX_split_join.sv:24:9
			wire [3:0] ipdom_tmask;
			// Trace: src/VX_split_join.sv:25:9
			wire [29:0] ipdom_pc;
			// Trace: src/VX_split_join.sv:26:9
			wire ipdom_idx;
			// Trace: src/VX_split_join.sv:27:9
			wire [33:0] ipdom_d0 = {split[37-:4] | split[33-:4], 30'sd0};
			// Trace: src/VX_split_join.sv:28:9
			wire [33:0] ipdom_d1 = {split[33-:4], split[29-:VX_gpu_pkg_PC_BITS]};
			// Trace: src/VX_split_join.sv:29:9
			wire sjoin_is_dvg = sjoin[1-:VX_gpu_pkg_DV_STACK_SIZEW] != ipdom_wr_ptr[wid * 2+:2];
			// Trace: src/VX_split_join.sv:30:9
			wire ipdom_push = split_valid && split[38];
			// Trace: src/VX_split_join.sv:31:9
			wire ipdom_pop = sjoin_valid && sjoin_is_dvg;
			// Trace: src/VX_split_join.sv:32:9
			VX_ipdom_stack #(
				.WIDTH(34),
				.DEPTH(VX_gpu_pkg_DV_STACK_SIZE)
			) ipdom_stack(
				.clk(clk),
				.reset(reset),
				.wid(wid),
				.d0(ipdom_d0),
				.d1(ipdom_d1),
				.push(ipdom_push),
				.pop(ipdom_pop),
				.rd_ptr(sjoin[1-:VX_gpu_pkg_DV_STACK_SIZEW]),
				.q_val({ipdom_tmask, ipdom_pc}),
				.q_idx(ipdom_idx),
				.wr_ptr(ipdom_wr_ptr),
				.empty(),
				.full()
			);
			// Trace: src/VX_split_join.sv:50:9
			VX_pipe_register #(
				.DATAW(39),
				.RESETW(1),
				.DEPTH(OUT_REG)
			) pipe_reg(
				.clk(clk),
				.reset(reset),
				.enable(1'b1),
				.data_in({sjoin_valid, wid, sjoin_is_dvg, ~ipdom_idx, ipdom_tmask, ipdom_pc}),
				.data_out({join_valid, join_wid, join_is_dvg, join_is_else, join_tmask, join_pc})
			);
			// Trace: src/VX_split_join.sv:61:9
			assign stack_ptr = ipdom_wr_ptr[stack_wid * 2+:2];
		end
	endgenerate
endmodule
// removed module with interface ports: VX_scoreboard
// removed module with interface ports: VX_wctl_unit
// removed module with interface ports: VX_alu_int
// removed interface: VX_issue_sched_if
// removed module with interface ports: VX_pe_switch
module VX_nz_iterator (
	clk,
	reset,
	valid_in,
	data_in,
	next,
	valid_out,
	data_out,
	pid,
	sop,
	eop
);
	// Trace: src/VX_nz_iterator.sv:2:13
	parameter DATAW = 8;
	// Trace: src/VX_nz_iterator.sv:3:13
	parameter KEYW = DATAW;
	// Trace: src/VX_nz_iterator.sv:4:13
	parameter N = 4;
	// Trace: src/VX_nz_iterator.sv:5:13
	parameter OUT_REG = 0;
	// Trace: src/VX_nz_iterator.sv:6:13
	parameter LPID_WIDTH = (N > 1 ? $clog2(N) : 1);
	// Trace: src/VX_nz_iterator.sv:8:5
	input wire clk;
	// Trace: src/VX_nz_iterator.sv:9:5
	input wire reset;
	// Trace: src/VX_nz_iterator.sv:10:5
	input wire valid_in;
	// Trace: src/VX_nz_iterator.sv:11:5
	input wire [(N * DATAW) - 1:0] data_in;
	// Trace: src/VX_nz_iterator.sv:12:5
	input wire next;
	// Trace: src/VX_nz_iterator.sv:13:5
	output wire valid_out;
	// Trace: src/VX_nz_iterator.sv:14:5
	output reg [DATAW - 1:0] data_out;
	// Trace: src/VX_nz_iterator.sv:15:5
	output reg [LPID_WIDTH - 1:0] pid;
	// Trace: src/VX_nz_iterator.sv:16:5
	output reg sop;
	// Trace: src/VX_nz_iterator.sv:17:5
	output reg eop;
	// Trace: src/VX_nz_iterator.sv:19:5
	function automatic signed [LPID_WIDTH - 1:0] sv2v_cast_54D48_signed;
		input reg signed [LPID_WIDTH - 1:0] inp;
		sv2v_cast_54D48_signed = inp;
	endfunction
	generate
		if (N > 1) begin : g_iterator
			// Trace: src/VX_nz_iterator.sv:20:9
			reg [N - 1:0] sent_mask_p;
			// Trace: src/VX_nz_iterator.sv:21:9
			wire [LPID_WIDTH - 1:0] start_p;
			wire [LPID_WIDTH - 1:0] end_p;
			// Trace: src/VX_nz_iterator.sv:22:9
			wire [N - 1:0] packet_valids;
			genvar _gv_i_152;
			for (_gv_i_152 = 0; _gv_i_152 < N; _gv_i_152 = _gv_i_152 + 1) begin : g_packet_valids
				localparam i = _gv_i_152;
				// Trace: src/VX_nz_iterator.sv:24:13
				assign packet_valids[i] = |data_in[(i * DATAW) + (KEYW - 1)-:KEYW];
			end
			// Trace: src/VX_nz_iterator.sv:26:9
			wire [(N * LPID_WIDTH) - 1:0] packet_ids;
			genvar _gv_i_153;
			for (_gv_i_153 = 0; _gv_i_153 < N; _gv_i_153 = _gv_i_153 + 1) begin : g_packet_ids
				localparam i = _gv_i_153;
				// Trace: src/VX_nz_iterator.sv:28:13
				assign packet_ids[i * LPID_WIDTH+:LPID_WIDTH] = sv2v_cast_54D48_signed(i);
			end
			// Trace: src/VX_nz_iterator.sv:30:9
			VX_find_first #(
				.N(N),
				.DATAW(LPID_WIDTH),
				.REVERSE(0)
			) find_first(
				.valid_in(packet_valids & ~sent_mask_p),
				.data_in(packet_ids),
				.data_out(start_p),
				.valid_out()
			);
			// Trace: src/VX_nz_iterator.sv:40:9
			VX_find_first #(
				.N(N),
				.DATAW(LPID_WIDTH),
				.REVERSE(1)
			) find_last(
				.valid_in(packet_valids),
				.data_in(packet_ids),
				.data_out(end_p),
				.valid_out()
			);
			// Trace: src/VX_nz_iterator.sv:50:9
			reg is_first_p;
			// Trace: src/VX_nz_iterator.sv:51:9
			wire is_last_p = start_p == end_p;
			// Trace: src/VX_nz_iterator.sv:52:9
			wire enable = valid_in && (~valid_out || next);
			// Trace: src/VX_nz_iterator.sv:53:9
			always @(posedge clk)
				// Trace: src/VX_nz_iterator.sv:54:13
				if (reset || (enable && (is_last_p || eop))) begin
					// Trace: src/VX_nz_iterator.sv:55:17
					sent_mask_p <= 1'sb0;
					// Trace: src/VX_nz_iterator.sv:56:17
					is_first_p <= 1;
				end
				else if (enable) begin
					// Trace: src/VX_nz_iterator.sv:58:17
					sent_mask_p[start_p] <= 1;
					// Trace: src/VX_nz_iterator.sv:59:17
					is_first_p <= 0;
				end
			// Trace: src/VX_nz_iterator.sv:62:9
			// rewrote reg-to-output bindings
			wire [((1 + DATAW) + LPID_WIDTH) + 2:1] sv2v_tmp_pipe_reg_data_out;
			always @(*) {valid_out, data_out, pid, sop, eop} = sv2v_tmp_pipe_reg_data_out;
			VX_pipe_register #(
				.DATAW(((1 + DATAW) + LPID_WIDTH) + 2),
				.RESETW(1),
				.DEPTH(OUT_REG)
			) pipe_reg(
				.clk(clk),
				.reset(reset || (enable && eop)),
				.enable(enable),
				.data_in({valid_in, data_in[start_p * DATAW+:DATAW], start_p, is_first_p, is_last_p}),
				.data_out(sv2v_tmp_pipe_reg_data_out)
			);
		end
		else begin : g_passthru
			// Trace: src/VX_nz_iterator.sv:74:9
			assign valid_out = valid_in;
			// Trace: src/VX_nz_iterator.sv:75:9
			wire [DATAW:1] sv2v_tmp_80DFB;
			assign sv2v_tmp_80DFB = data_in[0+:DATAW];
			always @(*) data_out = sv2v_tmp_80DFB;
			// Trace: src/VX_nz_iterator.sv:76:9
			wire [LPID_WIDTH:1] sv2v_tmp_1E98B;
			assign sv2v_tmp_1E98B = 0;
			always @(*) pid = sv2v_tmp_1E98B;
			// Trace: src/VX_nz_iterator.sv:77:9
			wire [1:1] sv2v_tmp_944DF;
			assign sv2v_tmp_944DF = 1;
			always @(*) sop = sv2v_tmp_944DF;
			// Trace: src/VX_nz_iterator.sv:78:9
			wire [1:1] sv2v_tmp_DEEF1;
			assign sv2v_tmp_DEEF1 = 1;
			always @(*) eop = sv2v_tmp_DEEF1;
		end
	endgenerate
endmodule
// removed module with interface ports: VX_csr_unit
module plru_decoder (
	way_idx,
	lru_data,
	lru_mask
);
	// removed import VX_gpu_pkg::*;
	// Trace: src/VX_cache_repl.sv:2:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_repl.sv:3:15
	parameter WAY_IDX_BITS = $clog2(NUM_WAYS);
	// Trace: src/VX_cache_repl.sv:4:15
	parameter WAY_IDX_WIDTH = (WAY_IDX_BITS > 0 ? WAY_IDX_BITS : 1);
	// Trace: src/VX_cache_repl.sv:6:5
	input wire [WAY_IDX_WIDTH - 1:0] way_idx;
	// Trace: src/VX_cache_repl.sv:7:5
	output wire [((NUM_WAYS - 1) > 0 ? NUM_WAYS - 1 : 1) - 1:0] lru_data;
	// Trace: src/VX_cache_repl.sv:8:5
	output wire [((NUM_WAYS - 1) > 0 ? NUM_WAYS - 1 : 1) - 1:0] lru_mask;
	// Trace: src/VX_cache_repl.sv:10:5
	generate
		if (NUM_WAYS > 1) begin : g_dec
			// Trace: src/VX_cache_repl.sv:11:9
			wire [((NUM_WAYS - 1) > 0 ? NUM_WAYS - 1 : 1) - 1:0] data;
			// Trace: src/VX_cache_repl.sv:12:9
			wire [((NUM_WAYS - 1) > 0 ? NUM_WAYS - 1 : 1) - 1:0] mask;
			genvar _gv_i_161;
			for (_gv_i_161 = 0; _gv_i_161 < (NUM_WAYS - 1); _gv_i_161 = _gv_i_161 + 1) begin : g_i
				localparam i = _gv_i_161;
				if (i == 0) begin : g_i_0
					// Trace: src/VX_cache_repl.sv:15:17
					assign mask[i] = 1'b1;
				end
				else if ((i % 2) == 1) begin : g_i_odd
					// Trace: src/VX_cache_repl.sv:17:17
					assign mask[i] = mask[(i - 1) / 2] & ~way_idx[(WAY_IDX_BITS - $clog2(i + 2)) + 1];
				end
				else begin : g_i_even
					// Trace: src/VX_cache_repl.sv:19:17
					assign mask[i] = mask[(i - 2) / 2] & way_idx[(WAY_IDX_BITS - $clog2(i + 2)) + 1];
				end
				// Trace: src/VX_cache_repl.sv:21:13
				assign data[i] = ~way_idx[WAY_IDX_BITS - $clog2(i + 2)];
			end
			// Trace: src/VX_cache_repl.sv:23:9
			assign lru_data = data;
			// Trace: src/VX_cache_repl.sv:24:9
			assign lru_mask = mask;
		end
		else begin : g_no_dec
			// Trace: src/VX_cache_repl.sv:26:9
			assign lru_data = 1'sb0;
			// Trace: src/VX_cache_repl.sv:27:9
			assign lru_mask = 1'sb0;
		end
	endgenerate
endmodule
module plru_encoder (
	lru_in,
	way_idx
);
	// Trace: src/VX_cache_repl.sv:31:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_repl.sv:32:15
	parameter WAY_IDX_BITS = $clog2(NUM_WAYS);
	// Trace: src/VX_cache_repl.sv:33:15
	parameter WAY_IDX_WIDTH = (WAY_IDX_BITS > 0 ? WAY_IDX_BITS : 1);
	// Trace: src/VX_cache_repl.sv:35:5
	input wire [((NUM_WAYS - 1) > 0 ? NUM_WAYS - 1 : 1) - 1:0] lru_in;
	// Trace: src/VX_cache_repl.sv:36:5
	output wire [WAY_IDX_WIDTH - 1:0] way_idx;
	// Trace: src/VX_cache_repl.sv:38:5
	generate
		if (NUM_WAYS > 1) begin : g_enc
			// Trace: src/VX_cache_repl.sv:39:9
			wire [WAY_IDX_BITS - 1:0] tmp;
			genvar _gv_i_162;
			for (_gv_i_162 = 0; _gv_i_162 < WAY_IDX_BITS; _gv_i_162 = _gv_i_162 + 1) begin : g_i
				localparam i = _gv_i_162;
				if (i == 0) begin : g_i_0
					// Trace: src/VX_cache_repl.sv:42:17
					assign tmp[WAY_IDX_WIDTH - 1] = lru_in[0];
				end
				else begin : g_i_n
					// Trace: src/VX_cache_repl.sv:44:17
					VX_mux #(.N(2 ** i)) mux(
						.data_in(lru_in[(2 ** i) - 1+:2 ** i]),
						.sel_in(tmp[WAY_IDX_BITS - 1-:i]),
						.data_out(tmp[(WAY_IDX_BITS - 1) - i])
					);
				end
			end
			// Trace: src/VX_cache_repl.sv:53:9
			assign way_idx = tmp;
		end
		else begin : g_no_enc
			// Trace: src/VX_cache_repl.sv:55:9
			assign way_idx = 1'sb0;
		end
	endgenerate
endmodule
module VX_cache_repl (
	clk,
	reset,
	stall,
	init,
	lookup_valid,
	lookup_hit,
	lookup_line,
	lookup_way,
	repl_valid,
	repl_line,
	repl_way
);
	// Trace: src/VX_cache_repl.sv:59:15
	parameter CACHE_SIZE = 1024;
	// Trace: src/VX_cache_repl.sv:60:15
	parameter LINE_SIZE = 64;
	// Trace: src/VX_cache_repl.sv:61:15
	parameter NUM_BANKS = 1;
	// Trace: src/VX_cache_repl.sv:62:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_repl.sv:63:15
	parameter REPL_POLICY = 1;
	// Trace: src/VX_cache_repl.sv:65:5
	input wire clk;
	// Trace: src/VX_cache_repl.sv:66:5
	input wire reset;
	// Trace: src/VX_cache_repl.sv:67:5
	input wire stall;
	// Trace: src/VX_cache_repl.sv:68:5
	input wire init;
	// Trace: src/VX_cache_repl.sv:69:5
	input wire lookup_valid;
	// Trace: src/VX_cache_repl.sv:70:5
	input wire lookup_hit;
	// Trace: src/VX_cache_repl.sv:71:5
	input wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] lookup_line;
	// Trace: src/VX_cache_repl.sv:72:5
	input wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] lookup_way;
	// Trace: src/VX_cache_repl.sv:73:5
	input wire repl_valid;
	// Trace: src/VX_cache_repl.sv:74:5
	input wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] repl_line;
	// Trace: src/VX_cache_repl.sv:75:5
	output wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] repl_way;
	// Trace: src/VX_cache_repl.sv:77:5
	localparam WAY_SEL_WIDTH = ($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1);
	// Trace: src/VX_cache_repl.sv:78:5
	generate
		if (NUM_WAYS > 1) begin : g_enable
			if (REPL_POLICY == 2) begin : g_plru
				// Trace: src/VX_cache_repl.sv:80:13
				localparam LRU_WIDTH = ((NUM_WAYS - 1) > 0 ? NUM_WAYS - 1 : 1);
				// Trace: src/VX_cache_repl.sv:81:13
				wire [LRU_WIDTH - 1:0] plru_rdata;
				// Trace: src/VX_cache_repl.sv:82:13
				wire [LRU_WIDTH - 1:0] plru_wdata;
				// Trace: src/VX_cache_repl.sv:83:13
				wire [LRU_WIDTH - 1:0] plru_wmask;
				// Trace: src/VX_cache_repl.sv:84:13
				localparam sv2v_uu_plru_store_WRENW = LRU_WIDTH;
				// removed localparam type sv2v_uu_plru_store_wren
				localparam [sv2v_uu_plru_store_WRENW - 1:0] sv2v_uu_plru_store_ext_wren_1 = 1'sb1;
				localparam sv2v_uu_plru_store_DATAW = LRU_WIDTH;
				// removed localparam type sv2v_uu_plru_store_wdata
				localparam [sv2v_uu_plru_store_DATAW - 1:0] sv2v_uu_plru_store_ext_wdata_0 = 1'sb0;
				VX_dp_ram #(
					.DATAW(LRU_WIDTH),
					.SIZE((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)),
					.WRENW(LRU_WIDTH),
					.RDW_MODE("R"),
					.RADDR_REG(1)
				) plru_store(
					.clk(clk),
					.reset(1'b0),
					.read(repl_valid),
					.write(init || (lookup_valid && lookup_hit)),
					.wren((init ? sv2v_uu_plru_store_ext_wren_1 : plru_wmask)),
					.waddr(lookup_line),
					.raddr(repl_line),
					.wdata((init ? sv2v_uu_plru_store_ext_wdata_0 : plru_wdata)),
					.rdata(plru_rdata)
				);
				// Trace: src/VX_cache_repl.sv:101:13
				plru_decoder #(.NUM_WAYS(NUM_WAYS)) plru_dec(
					.way_idx(lookup_way),
					.lru_data(plru_wdata),
					.lru_mask(plru_wmask)
				);
				// Trace: src/VX_cache_repl.sv:108:13
				plru_encoder #(.NUM_WAYS(NUM_WAYS)) plru_enc(
					.lru_in(plru_rdata),
					.way_idx(repl_way)
				);
			end
			else if (REPL_POLICY == 1) begin : g_fifo
				// Trace: src/VX_cache_repl.sv:115:13
				wire [WAY_SEL_WIDTH - 1:0] fifo_rdata;
				// Trace: src/VX_cache_repl.sv:116:13
				wire [WAY_SEL_WIDTH - 1:0] fifo_wdata = fifo_rdata + 1;
				// Trace: src/VX_cache_repl.sv:117:13
				localparam sv2v_uu_fifo_store_DATAW = WAY_SEL_WIDTH;
				// removed localparam type sv2v_uu_fifo_store_wdata
				localparam [sv2v_uu_fifo_store_DATAW - 1:0] sv2v_uu_fifo_store_ext_wdata_0 = 1'sb0;
				VX_sp_ram #(
					.DATAW(WAY_SEL_WIDTH),
					.SIZE((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)),
					.RDW_MODE("R"),
					.RADDR_REG(1)
				) fifo_store(
					.clk(clk),
					.reset(1'b0),
					.read(repl_valid),
					.write(init || repl_valid),
					.wren(1'b1),
					.addr(repl_line),
					.wdata((init ? sv2v_uu_fifo_store_ext_wdata_0 : fifo_wdata)),
					.rdata(fifo_rdata)
				);
				// Trace: src/VX_cache_repl.sv:132:13
				assign repl_way = fifo_rdata;
			end
			else begin : g_random
				// Trace: src/VX_cache_repl.sv:134:13
				reg [WAY_SEL_WIDTH - 1:0] victim_idx;
				// Trace: src/VX_cache_repl.sv:135:13
				always @(posedge clk)
					// Trace: src/VX_cache_repl.sv:136:17
					if (reset)
						// Trace: src/VX_cache_repl.sv:137:21
						victim_idx <= 0;
					else if (~stall)
						// Trace: src/VX_cache_repl.sv:139:21
						victim_idx <= victim_idx + 1;
				// Trace: src/VX_cache_repl.sv:142:13
				assign repl_way = victim_idx;
			end
		end
		else begin : g_disable
			// Trace: src/VX_cache_repl.sv:145:9
			assign repl_way = 1'b0;
		end
	endgenerate
endmodule
// removed interface: VX_result_if
// removed package "VX_trace_pkg"
module VX_popcount63 (
	data_in,
	data_out
);
	// Trace: src/VX_popcount.sv:2:5
	input wire [5:0] data_in;
	// Trace: src/VX_popcount.sv:3:5
	output wire [2:0] data_out;
	// Trace: src/VX_popcount.sv:5:5
	reg [2:0] sum;
	// Trace: src/VX_popcount.sv:6:5
	always @(*)
		// Trace: src/VX_popcount.sv:7:9
		case (data_in)
			6'd0:
				// Trace: src/VX_popcount.sv:8:16
				sum = 3'd0;
			6'd1:
				// Trace: src/VX_popcount.sv:8:34
				sum = 3'd1;
			6'd2:
				// Trace: src/VX_popcount.sv:8:52
				sum = 3'd1;
			6'd3:
				// Trace: src/VX_popcount.sv:8:70
				sum = 3'd2;
			6'd4:
				// Trace: src/VX_popcount.sv:9:16
				sum = 3'd1;
			6'd5:
				// Trace: src/VX_popcount.sv:9:34
				sum = 3'd2;
			6'd6:
				// Trace: src/VX_popcount.sv:9:52
				sum = 3'd2;
			6'd7:
				// Trace: src/VX_popcount.sv:9:70
				sum = 3'd3;
			6'd8:
				// Trace: src/VX_popcount.sv:10:16
				sum = 3'd1;
			6'd9:
				// Trace: src/VX_popcount.sv:10:34
				sum = 3'd2;
			6'd10:
				// Trace: src/VX_popcount.sv:10:52
				sum = 3'd2;
			6'd11:
				// Trace: src/VX_popcount.sv:10:70
				sum = 3'd3;
			6'd12:
				// Trace: src/VX_popcount.sv:11:16
				sum = 3'd2;
			6'd13:
				// Trace: src/VX_popcount.sv:11:34
				sum = 3'd3;
			6'd14:
				// Trace: src/VX_popcount.sv:11:52
				sum = 3'd3;
			6'd15:
				// Trace: src/VX_popcount.sv:11:70
				sum = 3'd4;
			6'd16:
				// Trace: src/VX_popcount.sv:12:16
				sum = 3'd1;
			6'd17:
				// Trace: src/VX_popcount.sv:12:34
				sum = 3'd2;
			6'd18:
				// Trace: src/VX_popcount.sv:12:52
				sum = 3'd2;
			6'd19:
				// Trace: src/VX_popcount.sv:12:70
				sum = 3'd3;
			6'd20:
				// Trace: src/VX_popcount.sv:13:16
				sum = 3'd2;
			6'd21:
				// Trace: src/VX_popcount.sv:13:34
				sum = 3'd3;
			6'd22:
				// Trace: src/VX_popcount.sv:13:52
				sum = 3'd3;
			6'd23:
				// Trace: src/VX_popcount.sv:13:70
				sum = 3'd4;
			6'd24:
				// Trace: src/VX_popcount.sv:14:16
				sum = 3'd2;
			6'd25:
				// Trace: src/VX_popcount.sv:14:34
				sum = 3'd3;
			6'd26:
				// Trace: src/VX_popcount.sv:14:52
				sum = 3'd3;
			6'd27:
				// Trace: src/VX_popcount.sv:14:70
				sum = 3'd4;
			6'd28:
				// Trace: src/VX_popcount.sv:15:16
				sum = 3'd3;
			6'd29:
				// Trace: src/VX_popcount.sv:15:34
				sum = 3'd4;
			6'd30:
				// Trace: src/VX_popcount.sv:15:52
				sum = 3'd4;
			6'd31:
				// Trace: src/VX_popcount.sv:15:70
				sum = 3'd5;
			6'd32:
				// Trace: src/VX_popcount.sv:16:16
				sum = 3'd1;
			6'd33:
				// Trace: src/VX_popcount.sv:16:34
				sum = 3'd2;
			6'd34:
				// Trace: src/VX_popcount.sv:16:52
				sum = 3'd2;
			6'd35:
				// Trace: src/VX_popcount.sv:16:70
				sum = 3'd3;
			6'd36:
				// Trace: src/VX_popcount.sv:17:16
				sum = 3'd2;
			6'd37:
				// Trace: src/VX_popcount.sv:17:34
				sum = 3'd3;
			6'd38:
				// Trace: src/VX_popcount.sv:17:52
				sum = 3'd3;
			6'd39:
				// Trace: src/VX_popcount.sv:17:70
				sum = 3'd4;
			6'd40:
				// Trace: src/VX_popcount.sv:18:16
				sum = 3'd2;
			6'd41:
				// Trace: src/VX_popcount.sv:18:34
				sum = 3'd3;
			6'd42:
				// Trace: src/VX_popcount.sv:18:52
				sum = 3'd3;
			6'd43:
				// Trace: src/VX_popcount.sv:18:70
				sum = 3'd4;
			6'd44:
				// Trace: src/VX_popcount.sv:19:16
				sum = 3'd3;
			6'd45:
				// Trace: src/VX_popcount.sv:19:34
				sum = 3'd4;
			6'd46:
				// Trace: src/VX_popcount.sv:19:52
				sum = 3'd4;
			6'd47:
				// Trace: src/VX_popcount.sv:19:70
				sum = 3'd5;
			6'd48:
				// Trace: src/VX_popcount.sv:20:16
				sum = 3'd2;
			6'd49:
				// Trace: src/VX_popcount.sv:20:34
				sum = 3'd3;
			6'd50:
				// Trace: src/VX_popcount.sv:20:52
				sum = 3'd3;
			6'd51:
				// Trace: src/VX_popcount.sv:20:70
				sum = 3'd4;
			6'd52:
				// Trace: src/VX_popcount.sv:21:16
				sum = 3'd3;
			6'd53:
				// Trace: src/VX_popcount.sv:21:34
				sum = 3'd4;
			6'd54:
				// Trace: src/VX_popcount.sv:21:52
				sum = 3'd4;
			6'd55:
				// Trace: src/VX_popcount.sv:21:70
				sum = 3'd5;
			6'd56:
				// Trace: src/VX_popcount.sv:22:16
				sum = 3'd3;
			6'd57:
				// Trace: src/VX_popcount.sv:22:34
				sum = 3'd4;
			6'd58:
				// Trace: src/VX_popcount.sv:22:52
				sum = 3'd4;
			6'd59:
				// Trace: src/VX_popcount.sv:22:70
				sum = 3'd5;
			6'd60:
				// Trace: src/VX_popcount.sv:23:16
				sum = 3'd4;
			6'd61:
				// Trace: src/VX_popcount.sv:23:34
				sum = 3'd5;
			6'd62:
				// Trace: src/VX_popcount.sv:23:52
				sum = 3'd5;
			6'd63:
				// Trace: src/VX_popcount.sv:23:70
				sum = 3'd6;
		endcase
	// Trace: src/VX_popcount.sv:26:5
	assign data_out = sum;
endmodule
module VX_popcount32 (
	data_in,
	data_out
);
	// Trace: src/VX_popcount.sv:29:5
	input wire [2:0] data_in;
	// Trace: src/VX_popcount.sv:30:5
	output wire [1:0] data_out;
	// Trace: src/VX_popcount.sv:32:5
	reg [1:0] sum;
	// Trace: src/VX_popcount.sv:33:5
	always @(*)
		// Trace: src/VX_popcount.sv:34:9
		case (data_in)
			3'd0:
				// Trace: src/VX_popcount.sv:35:15
				sum = 2'd0;
			3'd1:
				// Trace: src/VX_popcount.sv:35:33
				sum = 2'd1;
			3'd2:
				// Trace: src/VX_popcount.sv:35:51
				sum = 2'd1;
			3'd3:
				// Trace: src/VX_popcount.sv:35:69
				sum = 2'd2;
			3'd4:
				// Trace: src/VX_popcount.sv:36:15
				sum = 2'd1;
			3'd5:
				// Trace: src/VX_popcount.sv:36:33
				sum = 2'd2;
			3'd6:
				// Trace: src/VX_popcount.sv:36:51
				sum = 2'd2;
			3'd7:
				// Trace: src/VX_popcount.sv:36:69
				sum = 2'd3;
		endcase
	// Trace: src/VX_popcount.sv:39:5
	assign data_out = sum;
endmodule
module VX_sum33 (
	data_in1,
	data_in2,
	data_out
);
	// Trace: src/VX_popcount.sv:42:5
	input wire [2:0] data_in1;
	// Trace: src/VX_popcount.sv:43:5
	input wire [2:0] data_in2;
	// Trace: src/VX_popcount.sv:44:5
	output wire [3:0] data_out;
	// Trace: src/VX_popcount.sv:46:5
	reg [3:0] sum;
	// Trace: src/VX_popcount.sv:47:5
	always @(*)
		// Trace: src/VX_popcount.sv:48:9
		case ({data_in1, data_in2})
			6'd0:
				// Trace: src/VX_popcount.sv:49:16
				sum = 4'd0;
			6'd1:
				// Trace: src/VX_popcount.sv:49:34
				sum = 4'd1;
			6'd2:
				// Trace: src/VX_popcount.sv:49:52
				sum = 4'd2;
			6'd3:
				// Trace: src/VX_popcount.sv:49:70
				sum = 4'd3;
			6'd4:
				// Trace: src/VX_popcount.sv:50:16
				sum = 4'd4;
			6'd5:
				// Trace: src/VX_popcount.sv:50:34
				sum = 4'd5;
			6'd6:
				// Trace: src/VX_popcount.sv:50:52
				sum = 4'd6;
			6'd7:
				// Trace: src/VX_popcount.sv:50:70
				sum = 4'd7;
			6'd8:
				// Trace: src/VX_popcount.sv:51:16
				sum = 4'd1;
			6'd9:
				// Trace: src/VX_popcount.sv:51:34
				sum = 4'd2;
			6'd10:
				// Trace: src/VX_popcount.sv:51:52
				sum = 4'd3;
			6'd11:
				// Trace: src/VX_popcount.sv:51:70
				sum = 4'd4;
			6'd12:
				// Trace: src/VX_popcount.sv:52:16
				sum = 4'd5;
			6'd13:
				// Trace: src/VX_popcount.sv:52:34
				sum = 4'd6;
			6'd14:
				// Trace: src/VX_popcount.sv:52:52
				sum = 4'd7;
			6'd15:
				// Trace: src/VX_popcount.sv:52:70
				sum = 4'd8;
			6'd16:
				// Trace: src/VX_popcount.sv:53:16
				sum = 4'd2;
			6'd17:
				// Trace: src/VX_popcount.sv:53:34
				sum = 4'd3;
			6'd18:
				// Trace: src/VX_popcount.sv:53:52
				sum = 4'd4;
			6'd19:
				// Trace: src/VX_popcount.sv:53:70
				sum = 4'd5;
			6'd20:
				// Trace: src/VX_popcount.sv:54:16
				sum = 4'd6;
			6'd21:
				// Trace: src/VX_popcount.sv:54:34
				sum = 4'd7;
			6'd22:
				// Trace: src/VX_popcount.sv:54:52
				sum = 4'd8;
			6'd23:
				// Trace: src/VX_popcount.sv:54:70
				sum = 4'd9;
			6'd24:
				// Trace: src/VX_popcount.sv:55:16
				sum = 4'd3;
			6'd25:
				// Trace: src/VX_popcount.sv:55:34
				sum = 4'd4;
			6'd26:
				// Trace: src/VX_popcount.sv:55:52
				sum = 4'd5;
			6'd27:
				// Trace: src/VX_popcount.sv:55:70
				sum = 4'd6;
			6'd28:
				// Trace: src/VX_popcount.sv:56:16
				sum = 4'd7;
			6'd29:
				// Trace: src/VX_popcount.sv:56:34
				sum = 4'd8;
			6'd30:
				// Trace: src/VX_popcount.sv:56:52
				sum = 4'd9;
			6'd31:
				// Trace: src/VX_popcount.sv:56:70
				sum = 4'd10;
			6'd32:
				// Trace: src/VX_popcount.sv:57:16
				sum = 4'd4;
			6'd33:
				// Trace: src/VX_popcount.sv:57:34
				sum = 4'd5;
			6'd34:
				// Trace: src/VX_popcount.sv:57:52
				sum = 4'd6;
			6'd35:
				// Trace: src/VX_popcount.sv:57:70
				sum = 4'd7;
			6'd36:
				// Trace: src/VX_popcount.sv:58:16
				sum = 4'd8;
			6'd37:
				// Trace: src/VX_popcount.sv:58:34
				sum = 4'd9;
			6'd38:
				// Trace: src/VX_popcount.sv:58:52
				sum = 4'd10;
			6'd39:
				// Trace: src/VX_popcount.sv:58:70
				sum = 4'd11;
			6'd40:
				// Trace: src/VX_popcount.sv:59:16
				sum = 4'd5;
			6'd41:
				// Trace: src/VX_popcount.sv:59:34
				sum = 4'd6;
			6'd42:
				// Trace: src/VX_popcount.sv:59:52
				sum = 4'd7;
			6'd43:
				// Trace: src/VX_popcount.sv:59:70
				sum = 4'd8;
			6'd44:
				// Trace: src/VX_popcount.sv:60:16
				sum = 4'd9;
			6'd45:
				// Trace: src/VX_popcount.sv:60:34
				sum = 4'd10;
			6'd46:
				// Trace: src/VX_popcount.sv:60:52
				sum = 4'd11;
			6'd47:
				// Trace: src/VX_popcount.sv:60:70
				sum = 4'd12;
			6'd48:
				// Trace: src/VX_popcount.sv:61:16
				sum = 4'd6;
			6'd49:
				// Trace: src/VX_popcount.sv:61:34
				sum = 4'd7;
			6'd50:
				// Trace: src/VX_popcount.sv:61:52
				sum = 4'd8;
			6'd51:
				// Trace: src/VX_popcount.sv:61:70
				sum = 4'd9;
			6'd52:
				// Trace: src/VX_popcount.sv:62:16
				sum = 4'd10;
			6'd53:
				// Trace: src/VX_popcount.sv:62:34
				sum = 4'd11;
			6'd54:
				// Trace: src/VX_popcount.sv:62:52
				sum = 4'd12;
			6'd55:
				// Trace: src/VX_popcount.sv:62:70
				sum = 4'd13;
			6'd56:
				// Trace: src/VX_popcount.sv:63:16
				sum = 4'd7;
			6'd57:
				// Trace: src/VX_popcount.sv:63:34
				sum = 4'd8;
			6'd58:
				// Trace: src/VX_popcount.sv:63:52
				sum = 4'd9;
			6'd59:
				// Trace: src/VX_popcount.sv:63:70
				sum = 4'd10;
			6'd60:
				// Trace: src/VX_popcount.sv:64:16
				sum = 4'd11;
			6'd61:
				// Trace: src/VX_popcount.sv:64:34
				sum = 4'd12;
			6'd62:
				// Trace: src/VX_popcount.sv:64:52
				sum = 4'd13;
			6'd63:
				// Trace: src/VX_popcount.sv:64:70
				sum = 4'd14;
		endcase
	// Trace: src/VX_popcount.sv:67:5
	assign data_out = sum;
endmodule
module VX_popcount (
	data_in,
	data_out
);
	// Trace: src/VX_popcount.sv:70:15
	parameter MODEL = 1;
	// Trace: src/VX_popcount.sv:71:15
	parameter N = 1;
	// Trace: src/VX_popcount.sv:72:15
	parameter M = $clog2(N + 1);
	// Trace: src/VX_popcount.sv:74:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_popcount.sv:75:5
	output wire [M - 1:0] data_out;
	// Trace: src/VX_popcount.sv:77:5
	function automatic [M - 1:0] sv2v_cast_ABEB2;
		input reg [M - 1:0] inp;
		sv2v_cast_ABEB2 = inp;
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	generate
		if (N == 1) begin : g_passthru
			// Trace: src/VX_popcount.sv:78:9
			assign data_out = data_in;
		end
		else if (N <= 3) begin : g_popcount3
			// Trace: src/VX_popcount.sv:80:9
			reg [2:0] t_in;
			// Trace: src/VX_popcount.sv:81:9
			wire [1:0] t_out;
			// Trace: src/VX_popcount.sv:82:9
			always @(*) begin
				// Trace: src/VX_popcount.sv:83:13
				t_in = 1'sb0;
				// Trace: src/VX_popcount.sv:84:13
				t_in[N - 1:0] = data_in;
			end
			// Trace: src/VX_popcount.sv:86:9
			VX_popcount32 pc32(
				.data_in(t_in),
				.data_out(t_out)
			);
			// Trace: src/VX_popcount.sv:87:9
			assign data_out = t_out[M - 1:0];
		end
		else if (N <= 6) begin : g_popcount6
			// Trace: src/VX_popcount.sv:89:9
			reg [5:0] t_in;
			// Trace: src/VX_popcount.sv:90:9
			wire [2:0] t_out;
			// Trace: src/VX_popcount.sv:91:9
			always @(*) begin
				// Trace: src/VX_popcount.sv:92:13
				t_in = 1'sb0;
				// Trace: src/VX_popcount.sv:93:13
				t_in[N - 1:0] = data_in;
			end
			// Trace: src/VX_popcount.sv:95:9
			VX_popcount63 pc63(
				.data_in(t_in),
				.data_out(t_out)
			);
			// Trace: src/VX_popcount.sv:96:9
			assign data_out = t_out[M - 1:0];
		end
		else if (N <= 9) begin : g_popcount9
			// Trace: src/VX_popcount.sv:98:9
			reg [8:0] t_in;
			// Trace: src/VX_popcount.sv:99:9
			wire [4:0] t1_out;
			// Trace: src/VX_popcount.sv:100:9
			wire [3:0] t2_out;
			// Trace: src/VX_popcount.sv:101:9
			always @(*) begin
				// Trace: src/VX_popcount.sv:102:13
				t_in = 1'sb0;
				// Trace: src/VX_popcount.sv:103:13
				t_in[N - 1:0] = data_in;
			end
			// Trace: src/VX_popcount.sv:105:9
			VX_popcount63 pc63(
				.data_in(t_in[5:0]),
				.data_out(t1_out[2:0])
			);
			// Trace: src/VX_popcount.sv:106:9
			VX_popcount32 pc32(
				.data_in(t_in[8:6]),
				.data_out(t1_out[4:3])
			);
			// Trace: src/VX_popcount.sv:107:9
			VX_sum33 sum33(
				.data_in1(t1_out[2:0]),
				.data_in2({1'b0, t1_out[4:3]}),
				.data_out(t2_out)
			);
			// Trace: src/VX_popcount.sv:108:9
			assign data_out = t2_out[M - 1:0];
		end
		else if (N <= 12) begin : g_popcount12
			// Trace: src/VX_popcount.sv:110:9
			reg [11:0] t_in;
			// Trace: src/VX_popcount.sv:111:9
			wire [5:0] t1_out;
			// Trace: src/VX_popcount.sv:112:9
			wire [3:0] t2_out;
			// Trace: src/VX_popcount.sv:113:9
			always @(*) begin
				// Trace: src/VX_popcount.sv:114:13
				t_in = 1'sb0;
				// Trace: src/VX_popcount.sv:115:13
				t_in[N - 1:0] = data_in;
			end
			// Trace: src/VX_popcount.sv:117:9
			VX_popcount63 pc63a(
				.data_in(t_in[5:0]),
				.data_out(t1_out[2:0])
			);
			// Trace: src/VX_popcount.sv:118:9
			VX_popcount63 pc63b(
				.data_in(t_in[11:6]),
				.data_out(t1_out[5:3])
			);
			// Trace: src/VX_popcount.sv:119:9
			VX_sum33 sum33(
				.data_in1(t1_out[2:0]),
				.data_in2(t1_out[5:3]),
				.data_out(t2_out)
			);
			// Trace: src/VX_popcount.sv:120:9
			assign data_out = t2_out[M - 1:0];
		end
		else if (N <= 18) begin : g_popcount18
			// Trace: src/VX_popcount.sv:122:9
			reg [17:0] t_in;
			// Trace: src/VX_popcount.sv:123:9
			wire [8:0] t1_out;
			// Trace: src/VX_popcount.sv:124:9
			wire [5:0] t2_out;
			// Trace: src/VX_popcount.sv:125:9
			always @(*) begin
				// Trace: src/VX_popcount.sv:126:13
				t_in = 1'sb0;
				// Trace: src/VX_popcount.sv:127:13
				t_in[N - 1:0] = data_in;
			end
			// Trace: src/VX_popcount.sv:129:9
			VX_popcount63 pc63a(
				.data_in(t_in[5:0]),
				.data_out(t1_out[2:0])
			);
			// Trace: src/VX_popcount.sv:130:9
			VX_popcount63 pc63b(
				.data_in(t_in[11:6]),
				.data_out(t1_out[5:3])
			);
			// Trace: src/VX_popcount.sv:131:9
			VX_popcount63 pc63c(
				.data_in(t_in[17:12]),
				.data_out(t1_out[8:6])
			);
			// Trace: src/VX_popcount.sv:132:9
			VX_popcount32 pc32a(
				.data_in({t1_out[0], t1_out[3], t1_out[6]}),
				.data_out(t2_out[1:0])
			);
			// Trace: src/VX_popcount.sv:133:9
			VX_popcount32 pc32b(
				.data_in({t1_out[1], t1_out[4], t1_out[7]}),
				.data_out(t2_out[3:2])
			);
			// Trace: src/VX_popcount.sv:134:9
			VX_popcount32 pc32c(
				.data_in({t1_out[2], t1_out[5], t1_out[8]}),
				.data_out(t2_out[5:4])
			);
			// Trace: src/VX_popcount.sv:135:9
			assign data_out = ({2'b00, t2_out[1:0]} + {1'b0, t2_out[3:2], 1'b0}) + {t2_out[5:4], 2'b00};
		end
		else if (MODEL == 1) begin : g_model1
			// Trace: src/VX_popcount.sv:137:9
			localparam PN = 1 << $clog2(N);
			// Trace: src/VX_popcount.sv:138:9
			localparam LOGPN = $clog2(PN);
			// Trace: src/VX_popcount.sv:139:9
			wire [M - 1:0] tmp [LOGPN - 1:0][PN - 1:0];
			genvar _gv_j_18;
			for (_gv_j_18 = 0; _gv_j_18 < LOGPN; _gv_j_18 = _gv_j_18 + 1) begin : genblk1
				localparam j = _gv_j_18;
				// Trace: src/VX_popcount.sv:141:13
				localparam D = j + 1;
				// Trace: src/VX_popcount.sv:142:13
				localparam Q = (D < LOGPN ? D + 1 : M);
				genvar _gv_i_171;
				for (_gv_i_171 = 0; _gv_i_171 < (1 << ((LOGPN - j) - 1)); _gv_i_171 = _gv_i_171 + 1) begin : genblk1
					localparam i = _gv_i_171;
					// Trace: src/VX_popcount.sv:144:17
					localparam l = i * 2;
					// Trace: src/VX_popcount.sv:145:17
					localparam r = (i * 2) + 1;
					// Trace: src/VX_popcount.sv:146:17
					wire [Q - 1:0] res;
					if (j == 0) begin : genblk1
						if (r < N) begin : genblk1
							// Trace: src/VX_popcount.sv:149:25
							assign res = data_in[l] + data_in[r];
						end
						else if (l < N) begin : genblk1
							// Trace: src/VX_popcount.sv:151:25
							assign res = sv2v_cast_2(data_in[l]);
						end
						else begin : genblk1
							// Trace: src/VX_popcount.sv:153:25
							assign res = 2'b00;
						end
					end
					else begin : genblk1
						// Trace: src/VX_popcount.sv:156:21
						function automatic [D - 1:0] sv2v_cast_AC9B9;
							input reg [D - 1:0] inp;
							sv2v_cast_AC9B9 = inp;
						endfunction
						assign res = sv2v_cast_AC9B9(tmp[j - 1][l]) + sv2v_cast_AC9B9(tmp[j - 1][r]);
					end
					// Trace: src/VX_popcount.sv:158:17
					assign tmp[j][i] = sv2v_cast_ABEB2(res);
				end
			end
			// Trace: src/VX_popcount.sv:161:9
			assign data_out = tmp[LOGPN - 1][0];
		end
		else begin : g_model2
			// Trace: src/VX_popcount.sv:163:9
			reg [M - 1:0] cnt_w;
			// Trace: src/VX_popcount.sv:164:9
			always @(*) begin
				// Trace: src/VX_popcount.sv:165:13
				cnt_w = 1'sb0;
				// Trace: src/VX_popcount.sv:166:13
				begin : sv2v_autoblock_1
					// Trace: src/VX_popcount.sv:166:18
					integer i;
					// Trace: src/VX_popcount.sv:166:18
					for (i = 0; i < N; i = i + 1)
						begin
							// Trace: src/VX_popcount.sv:167:17
							cnt_w = cnt_w + sv2v_cast_ABEB2(data_in[i]);
						end
				end
			end
			// Trace: src/VX_popcount.sv:170:9
			assign data_out = cnt_w;
		end
	endgenerate
endmodule
// removed interface: VX_warp_ctl_if
// removed module with interface ports: VX_lsu_adapter
// removed module with interface ports: VX_socket
// removed module with interface ports: VX_gbar_arb
// removed module with interface ports: VX_mem_arb
// removed interface: VX_sched_csr_if
// removed interface: VX_execute_if
// removed interface: VX_operands_if
// removed module with interface ports: VX_lsu_unit
// removed module with interface ports: VX_cache_cluster
module VX_stream_unpack (
	clk,
	reset,
	valid_in,
	mask_in,
	data_in,
	tag_in,
	ready_in,
	valid_out,
	data_out,
	tag_out,
	ready_out
);
	// Trace: src/VX_stream_unpack.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_stream_unpack.sv:3:15
	parameter DATA_WIDTH = 1;
	// Trace: src/VX_stream_unpack.sv:4:15
	parameter TAG_WIDTH = 1;
	// Trace: src/VX_stream_unpack.sv:5:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_stream_unpack.sv:7:5
	input wire clk;
	// Trace: src/VX_stream_unpack.sv:8:5
	input wire reset;
	// Trace: src/VX_stream_unpack.sv:9:5
	input wire valid_in;
	// Trace: src/VX_stream_unpack.sv:10:5
	input wire [NUM_REQS - 1:0] mask_in;
	// Trace: src/VX_stream_unpack.sv:11:5
	input wire [(NUM_REQS * DATA_WIDTH) - 1:0] data_in;
	// Trace: src/VX_stream_unpack.sv:12:5
	input wire [TAG_WIDTH - 1:0] tag_in;
	// Trace: src/VX_stream_unpack.sv:13:5
	output wire ready_in;
	// Trace: src/VX_stream_unpack.sv:14:5
	output wire [NUM_REQS - 1:0] valid_out;
	// Trace: src/VX_stream_unpack.sv:15:5
	output wire [(NUM_REQS * DATA_WIDTH) - 1:0] data_out;
	// Trace: src/VX_stream_unpack.sv:16:5
	output wire [(NUM_REQS * TAG_WIDTH) - 1:0] tag_out;
	// Trace: src/VX_stream_unpack.sv:17:5
	input wire [NUM_REQS - 1:0] ready_out;
	// Trace: src/VX_stream_unpack.sv:19:5
	generate
		if (NUM_REQS > 1) begin : g_unpack
			// Trace: src/VX_stream_unpack.sv:20:9
			reg [NUM_REQS - 1:0] rem_mask_r;
			// Trace: src/VX_stream_unpack.sv:21:9
			wire [NUM_REQS - 1:0] ready_out_w;
			// Trace: src/VX_stream_unpack.sv:22:9
			wire [NUM_REQS - 1:0] rem_mask_n = rem_mask_r & ~ready_out_w;
			// Trace: src/VX_stream_unpack.sv:23:9
			wire sent_all = ~(|(mask_in & rem_mask_n));
			// Trace: src/VX_stream_unpack.sv:24:9
			always @(posedge clk)
				// Trace: src/VX_stream_unpack.sv:25:13
				if (reset)
					// Trace: src/VX_stream_unpack.sv:26:17
					rem_mask_r <= 1'sb1;
				else
					// Trace: src/VX_stream_unpack.sv:28:17
					if (valid_in)
						// Trace: src/VX_stream_unpack.sv:29:21
						rem_mask_r <= (sent_all ? {NUM_REQS {1'sb1}} : rem_mask_n);
			// Trace: src/VX_stream_unpack.sv:33:9
			assign ready_in = sent_all;
			genvar _gv_i_194;
			for (_gv_i_194 = 0; _gv_i_194 < NUM_REQS; _gv_i_194 = _gv_i_194 + 1) begin : g_outbuf
				localparam i = _gv_i_194;
				// Trace: src/VX_stream_unpack.sv:35:13
				VX_elastic_buffer #(
					.DATAW(DATA_WIDTH + TAG_WIDTH),
					.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
					.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
				) out_buf(
					.clk(clk),
					.reset(reset),
					.valid_in((valid_in && mask_in[i]) && rem_mask_r[i]),
					.ready_in(ready_out_w[i]),
					.data_in({data_in[i * DATA_WIDTH+:DATA_WIDTH], tag_in}),
					.data_out({data_out[i * DATA_WIDTH+:DATA_WIDTH], tag_out[i * TAG_WIDTH+:TAG_WIDTH]}),
					.valid_out(valid_out[i]),
					.ready_out(ready_out[i])
				);
			end
		end
		else begin : g_passthru
			// Trace: src/VX_stream_unpack.sv:51:9
			assign valid_out = valid_in;
			// Trace: src/VX_stream_unpack.sv:52:9
			assign data_out = data_in;
			// Trace: src/VX_stream_unpack.sv:53:9
			assign tag_out = tag_in;
			// Trace: src/VX_stream_unpack.sv:54:9
			assign ready_in = ready_out;
		end
	endgenerate
endmodule
module VX_cache_bank (
	clk,
	reset,
	core_req_valid,
	core_req_addr,
	core_req_rw,
	core_req_wsel,
	core_req_byteen,
	core_req_data,
	core_req_tag,
	core_req_idx,
	core_req_flags,
	core_req_ready,
	core_rsp_valid,
	core_rsp_data,
	core_rsp_tag,
	core_rsp_idx,
	core_rsp_ready,
	mem_req_valid,
	mem_req_addr,
	mem_req_rw,
	mem_req_byteen,
	mem_req_data,
	mem_req_tag,
	mem_req_flags,
	mem_req_ready,
	mem_rsp_valid,
	mem_rsp_data,
	mem_rsp_tag,
	mem_rsp_ready,
	flush_begin,
	flush_uuid,
	flush_end
);
	// removed import VX_gpu_pkg::*;
	// Trace: src/VX_cache_bank.sv:2:15
	parameter INSTANCE_ID = "";
	// Trace: src/VX_cache_bank.sv:3:15
	parameter BANK_ID = 0;
	// Trace: src/VX_cache_bank.sv:4:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_cache_bank.sv:5:15
	parameter CACHE_SIZE = 1024;
	// Trace: src/VX_cache_bank.sv:6:15
	parameter LINE_SIZE = 16;
	// Trace: src/VX_cache_bank.sv:7:15
	parameter NUM_BANKS = 1;
	// Trace: src/VX_cache_bank.sv:8:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_bank.sv:9:15
	parameter WORD_SIZE = 4;
	// Trace: src/VX_cache_bank.sv:10:15
	parameter CRSQ_SIZE = 1;
	// Trace: src/VX_cache_bank.sv:11:15
	parameter MSHR_SIZE = 1;
	// Trace: src/VX_cache_bank.sv:12:15
	parameter MREQ_SIZE = 1;
	// Trace: src/VX_cache_bank.sv:13:15
	parameter WRITE_ENABLE = 1;
	// Trace: src/VX_cache_bank.sv:14:15
	parameter WRITEBACK = 0;
	// Trace: src/VX_cache_bank.sv:15:15
	parameter DIRTY_BYTES = 0;
	// Trace: src/VX_cache_bank.sv:16:15
	parameter REPL_POLICY = 1;
	// Trace: src/VX_cache_bank.sv:17:15
	localparam VX_gpu_pkg_UUID_WIDTH = 1;
	parameter TAG_WIDTH = 2;
	// Trace: src/VX_cache_bank.sv:18:15
	parameter CORE_OUT_REG = 0;
	// Trace: src/VX_cache_bank.sv:19:15
	parameter MEM_OUT_REG = 0;
	// Trace: src/VX_cache_bank.sv:20:15
	parameter MSHR_ADDR_WIDTH = (MSHR_SIZE > 1 ? $clog2(MSHR_SIZE) : 1);
	// Trace: src/VX_cache_bank.sv:21:15
	parameter MEM_TAG_WIDTH = VX_gpu_pkg_UUID_WIDTH + MSHR_ADDR_WIDTH;
	// Trace: src/VX_cache_bank.sv:22:15
	parameter REQ_SEL_WIDTH = ($clog2(NUM_REQS) > 0 ? $clog2(NUM_REQS) : 1);
	// Trace: src/VX_cache_bank.sv:23:15
	parameter WORD_SEL_WIDTH = ($clog2(LINE_SIZE / WORD_SIZE) > 0 ? $clog2(LINE_SIZE / WORD_SIZE) : 1);
	// Trace: src/VX_cache_bank.sv:25:5
	input wire clk;
	// Trace: src/VX_cache_bank.sv:26:5
	input wire reset;
	// Trace: src/VX_cache_bank.sv:27:5
	input wire core_req_valid;
	// Trace: src/VX_cache_bank.sv:28:5
	input wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] core_req_addr;
	// Trace: src/VX_cache_bank.sv:29:5
	input wire core_req_rw;
	// Trace: src/VX_cache_bank.sv:30:5
	input wire [WORD_SEL_WIDTH - 1:0] core_req_wsel;
	// Trace: src/VX_cache_bank.sv:31:5
	input wire [WORD_SIZE - 1:0] core_req_byteen;
	// Trace: src/VX_cache_bank.sv:32:5
	input wire [(8 * WORD_SIZE) - 1:0] core_req_data;
	// Trace: src/VX_cache_bank.sv:33:5
	input wire [TAG_WIDTH - 1:0] core_req_tag;
	// Trace: src/VX_cache_bank.sv:34:5
	input wire [REQ_SEL_WIDTH - 1:0] core_req_idx;
	// Trace: src/VX_cache_bank.sv:35:5
	localparam VX_gpu_pkg_MEM_REQ_FLAG_LOCAL = 2;
	localparam VX_gpu_pkg_MEM_FLAGS_WIDTH = 3;
	input wire [2:0] core_req_flags;
	// Trace: src/VX_cache_bank.sv:36:5
	output wire core_req_ready;
	// Trace: src/VX_cache_bank.sv:37:5
	output wire core_rsp_valid;
	// Trace: src/VX_cache_bank.sv:38:5
	output wire [(8 * WORD_SIZE) - 1:0] core_rsp_data;
	// Trace: src/VX_cache_bank.sv:39:5
	output wire [TAG_WIDTH - 1:0] core_rsp_tag;
	// Trace: src/VX_cache_bank.sv:40:5
	output wire [REQ_SEL_WIDTH - 1:0] core_rsp_idx;
	// Trace: src/VX_cache_bank.sv:41:5
	input wire core_rsp_ready;
	// Trace: src/VX_cache_bank.sv:42:5
	output wire mem_req_valid;
	// Trace: src/VX_cache_bank.sv:43:5
	output wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] mem_req_addr;
	// Trace: src/VX_cache_bank.sv:44:5
	output wire mem_req_rw;
	// Trace: src/VX_cache_bank.sv:45:5
	output wire [LINE_SIZE - 1:0] mem_req_byteen;
	// Trace: src/VX_cache_bank.sv:46:5
	output wire [(8 * LINE_SIZE) - 1:0] mem_req_data;
	// Trace: src/VX_cache_bank.sv:47:5
	output wire [MEM_TAG_WIDTH - 1:0] mem_req_tag;
	// Trace: src/VX_cache_bank.sv:48:5
	output wire [2:0] mem_req_flags;
	// Trace: src/VX_cache_bank.sv:49:5
	input wire mem_req_ready;
	// Trace: src/VX_cache_bank.sv:50:5
	input wire mem_rsp_valid;
	// Trace: src/VX_cache_bank.sv:51:5
	input wire [(8 * LINE_SIZE) - 1:0] mem_rsp_data;
	// Trace: src/VX_cache_bank.sv:52:5
	input wire [MEM_TAG_WIDTH - 1:0] mem_rsp_tag;
	// Trace: src/VX_cache_bank.sv:53:5
	output wire mem_rsp_ready;
	// Trace: src/VX_cache_bank.sv:54:5
	input wire flush_begin;
	// Trace: src/VX_cache_bank.sv:55:5
	input wire [0:0] flush_uuid;
	// Trace: src/VX_cache_bank.sv:56:5
	output wire flush_end;
	// Trace: src/VX_cache_bank.sv:58:5
	localparam PIPELINE_STAGES = 2;
	// Trace: src/VX_cache_bank.sv:59:5
	wire [0:0] req_uuid_sel;
	wire [0:0] req_uuid_st0;
	wire [0:0] req_uuid_st1;
	// Trace: src/VX_cache_bank.sv:60:5
	wire crsp_queue_stall;
	// Trace: src/VX_cache_bank.sv:61:5
	wire mshr_alm_full;
	// Trace: src/VX_cache_bank.sv:62:5
	wire mreq_queue_empty;
	// Trace: src/VX_cache_bank.sv:63:5
	wire mreq_queue_alm_full;
	// Trace: src/VX_cache_bank.sv:64:5
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] mem_rsp_addr;
	// Trace: src/VX_cache_bank.sv:65:5
	wire replay_valid;
	// Trace: src/VX_cache_bank.sv:66:5
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] replay_addr;
	// Trace: src/VX_cache_bank.sv:67:5
	wire replay_rw;
	// Trace: src/VX_cache_bank.sv:68:5
	wire [WORD_SEL_WIDTH - 1:0] replay_wsel;
	// Trace: src/VX_cache_bank.sv:69:5
	wire [WORD_SIZE - 1:0] replay_byteen;
	// Trace: src/VX_cache_bank.sv:70:5
	wire [(8 * WORD_SIZE) - 1:0] replay_data;
	// Trace: src/VX_cache_bank.sv:71:5
	wire [TAG_WIDTH - 1:0] replay_tag;
	// Trace: src/VX_cache_bank.sv:72:5
	wire [REQ_SEL_WIDTH - 1:0] replay_idx;
	// Trace: src/VX_cache_bank.sv:73:5
	wire [MSHR_ADDR_WIDTH - 1:0] replay_id;
	// Trace: src/VX_cache_bank.sv:74:5
	wire replay_ready;
	// Trace: src/VX_cache_bank.sv:75:5
	wire valid_sel;
	wire valid_st0;
	wire valid_st1;
	// Trace: src/VX_cache_bank.sv:76:5
	wire is_init_st0;
	// Trace: src/VX_cache_bank.sv:77:5
	wire is_creq_st0;
	wire is_creq_st1;
	// Trace: src/VX_cache_bank.sv:78:5
	wire is_fill_st0;
	wire is_fill_st1;
	// Trace: src/VX_cache_bank.sv:79:5
	wire is_flush_st0;
	wire is_flush_st1;
	// Trace: src/VX_cache_bank.sv:80:5
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] flush_way_st0;
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] evict_way_st0;
	// Trace: src/VX_cache_bank.sv:81:5
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] way_idx_st0;
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] way_idx_st1;
	// Trace: src/VX_cache_bank.sv:82:5
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] addr_sel;
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] addr_st0;
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] addr_st1;
	// Trace: src/VX_cache_bank.sv:83:5
	wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] line_idx_sel;
	wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] line_idx_st0;
	wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] line_idx_st1;
	// Trace: src/VX_cache_bank.sv:84:5
	wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) - 1:0] line_tag_st0;
	wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) - 1:0] line_tag_st1;
	// Trace: src/VX_cache_bank.sv:85:5
	wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) - 1:0] evict_tag_st0;
	wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) - 1:0] evict_tag_st1;
	// Trace: src/VX_cache_bank.sv:86:5
	wire rw_sel;
	wire rw_st0;
	wire rw_st1;
	// Trace: src/VX_cache_bank.sv:87:5
	wire [WORD_SEL_WIDTH - 1:0] word_idx_sel;
	wire [WORD_SEL_WIDTH - 1:0] word_idx_st0;
	wire [WORD_SEL_WIDTH - 1:0] word_idx_st1;
	// Trace: src/VX_cache_bank.sv:88:5
	wire [WORD_SIZE - 1:0] byteen_sel;
	wire [WORD_SIZE - 1:0] byteen_st0;
	wire [WORD_SIZE - 1:0] byteen_st1;
	// Trace: src/VX_cache_bank.sv:89:5
	wire [REQ_SEL_WIDTH - 1:0] req_idx_sel;
	wire [REQ_SEL_WIDTH - 1:0] req_idx_st0;
	wire [REQ_SEL_WIDTH - 1:0] req_idx_st1;
	// Trace: src/VX_cache_bank.sv:90:5
	wire [TAG_WIDTH - 1:0] tag_sel;
	wire [TAG_WIDTH - 1:0] tag_st0;
	wire [TAG_WIDTH - 1:0] tag_st1;
	// Trace: src/VX_cache_bank.sv:91:5
	wire [(8 * WORD_SIZE) - 1:0] write_word_st0;
	wire [(8 * WORD_SIZE) - 1:0] write_word_st1;
	// Trace: src/VX_cache_bank.sv:92:5
	wire [(8 * LINE_SIZE) - 1:0] data_sel;
	wire [(8 * LINE_SIZE) - 1:0] data_st0;
	wire [(8 * LINE_SIZE) - 1:0] data_st1;
	// Trace: src/VX_cache_bank.sv:93:5
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_id_st0;
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_id_st1;
	// Trace: src/VX_cache_bank.sv:94:5
	wire [MSHR_ADDR_WIDTH - 1:0] replay_id_st0;
	// Trace: src/VX_cache_bank.sv:95:5
	wire is_dirty_st0;
	wire is_dirty_st1;
	// Trace: src/VX_cache_bank.sv:96:5
	wire is_replay_st0;
	wire is_replay_st1;
	// Trace: src/VX_cache_bank.sv:97:5
	wire is_hit_st0;
	wire is_hit_st1;
	// Trace: src/VX_cache_bank.sv:98:5
	wire [2:0] flags_sel;
	wire [2:0] flags_st0;
	wire [2:0] flags_st1;
	// Trace: src/VX_cache_bank.sv:99:5
	wire mshr_pending_st0;
	wire mshr_pending_st1;
	// Trace: src/VX_cache_bank.sv:100:5
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_previd_st0;
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_previd_st1;
	// Trace: src/VX_cache_bank.sv:101:5
	wire mshr_empty;
	// Trace: src/VX_cache_bank.sv:102:5
	wire flush_valid;
	// Trace: src/VX_cache_bank.sv:103:5
	wire init_valid;
	// Trace: src/VX_cache_bank.sv:104:5
	wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] flush_sel;
	// Trace: src/VX_cache_bank.sv:105:5
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] flush_way;
	// Trace: src/VX_cache_bank.sv:106:5
	wire flush_ready;
	// Trace: src/VX_cache_bank.sv:107:5
	wire no_pending_req = (~valid_st0 && ~valid_st1) && mreq_queue_empty;
	// Trace: src/VX_cache_bank.sv:108:5
	VX_cache_flush #(
		.BANK_ID(BANK_ID),
		.CACHE_SIZE(CACHE_SIZE),
		.LINE_SIZE(LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.NUM_WAYS(NUM_WAYS),
		.WRITEBACK(WRITEBACK)
	) cache_flush(
		.clk(clk),
		.reset(reset),
		.flush_begin(flush_begin),
		.flush_end(flush_end),
		.flush_init(init_valid),
		.flush_valid(flush_valid),
		.flush_line(flush_sel),
		.flush_way(flush_way),
		.flush_ready(flush_ready),
		.mshr_empty(mshr_empty),
		.bank_empty(no_pending_req)
	);
	// Trace: src/VX_cache_bank.sv:128:5
	wire pipe_stall = crsp_queue_stall;
	// Trace: src/VX_cache_bank.sv:129:5
	wire replay_grant = ~init_valid;
	// Trace: src/VX_cache_bank.sv:130:5
	wire replay_enable = replay_grant && replay_valid;
	// Trace: src/VX_cache_bank.sv:131:5
	wire fill_grant = ~init_valid && ~replay_enable;
	// Trace: src/VX_cache_bank.sv:132:5
	wire fill_enable = fill_grant && mem_rsp_valid;
	// Trace: src/VX_cache_bank.sv:133:5
	wire flush_grant = (~init_valid && ~replay_enable) && ~fill_enable;
	// Trace: src/VX_cache_bank.sv:134:5
	wire flush_enable = flush_grant && flush_valid;
	// Trace: src/VX_cache_bank.sv:135:5
	wire creq_grant = ((~init_valid && ~replay_enable) && ~fill_enable) && ~flush_enable;
	// Trace: src/VX_cache_bank.sv:136:5
	wire creq_enable = creq_grant && core_req_valid;
	// Trace: src/VX_cache_bank.sv:137:5
	assign replay_ready = (replay_grant && ~((!WRITEBACK && replay_rw) && mreq_queue_alm_full)) && ~pipe_stall;
	// Trace: src/VX_cache_bank.sv:140:5
	assign mem_rsp_ready = (fill_grant && ~(WRITEBACK && mreq_queue_alm_full)) && ~pipe_stall;
	// Trace: src/VX_cache_bank.sv:143:5
	assign flush_ready = (flush_grant && ~(WRITEBACK && mreq_queue_alm_full)) && ~pipe_stall;
	// Trace: src/VX_cache_bank.sv:146:5
	assign core_req_ready = ((creq_grant && ~mreq_queue_alm_full) && ~mshr_alm_full) && ~pipe_stall;
	// Trace: src/VX_cache_bank.sv:150:5
	wire init_fire = init_valid;
	// Trace: src/VX_cache_bank.sv:151:5
	wire replay_fire = replay_valid && replay_ready;
	// Trace: src/VX_cache_bank.sv:152:5
	wire mem_rsp_fire = mem_rsp_valid && mem_rsp_ready;
	// Trace: src/VX_cache_bank.sv:153:5
	wire flush_fire = flush_valid && flush_ready;
	// Trace: src/VX_cache_bank.sv:154:5
	wire core_req_fire = core_req_valid && core_req_ready;
	// Trace: src/VX_cache_bank.sv:155:5
	wire [MSHR_ADDR_WIDTH - 1:0] mem_rsp_id = mem_rsp_tag[MSHR_ADDR_WIDTH - 1:0];
	// Trace: src/VX_cache_bank.sv:156:5
	wire [TAG_WIDTH - 1:0] mem_rsp_tag_s;
	// Trace: src/VX_cache_bank.sv:157:5
	function automatic [(TAG_WIDTH - MEM_TAG_WIDTH) - 1:0] sv2v_cast_E6004;
		input reg [(TAG_WIDTH - MEM_TAG_WIDTH) - 1:0] inp;
		sv2v_cast_E6004 = inp;
	endfunction
	generate
		if (TAG_WIDTH > MEM_TAG_WIDTH) begin : g_mem_rsp_tag_s_pad
			// Trace: src/VX_cache_bank.sv:158:9
			assign mem_rsp_tag_s = {mem_rsp_tag, sv2v_cast_E6004(1'b0)};
		end
		else begin : g_mem_rsp_tag_s_cut
			// Trace: src/VX_cache_bank.sv:160:9
			assign mem_rsp_tag_s = mem_rsp_tag[MEM_TAG_WIDTH - 1-:TAG_WIDTH];
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:162:5
	wire [TAG_WIDTH - 1:0] flush_tag;
	// Trace: src/VX_cache_bank.sv:163:5
	function automatic [((TAG_WIDTH - 2) >= 0 ? TAG_WIDTH - 1 : 3 - TAG_WIDTH) - 1:0] sv2v_cast_756E4;
		input reg [((TAG_WIDTH - 2) >= 0 ? TAG_WIDTH - 1 : 3 - TAG_WIDTH) - 1:0] inp;
		sv2v_cast_756E4 = inp;
	endfunction
	generate
		if (1) begin : g_flush_tag_uuid
			// Trace: src/VX_cache_bank.sv:164:9
			assign flush_tag = {flush_uuid, sv2v_cast_756E4(1'b0)};
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:168:5
	assign valid_sel = (((init_fire || replay_fire) || mem_rsp_fire) || flush_fire) || core_req_fire;
	// Trace: src/VX_cache_bank.sv:169:5
	assign rw_sel = (replay_valid ? replay_rw : core_req_rw);
	// Trace: src/VX_cache_bank.sv:170:5
	assign byteen_sel = (replay_valid ? replay_byteen : core_req_byteen);
	// Trace: src/VX_cache_bank.sv:171:5
	function automatic [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] sv2v_cast_9CD28;
		input reg [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] inp;
		sv2v_cast_9CD28 = inp;
	endfunction
	assign addr_sel = (init_valid | flush_valid ? sv2v_cast_9CD28(flush_sel) : (replay_valid ? replay_addr : (mem_rsp_valid ? mem_rsp_addr : core_req_addr)));
	// Trace: src/VX_cache_bank.sv:173:5
	assign word_idx_sel = (replay_valid ? replay_wsel : core_req_wsel);
	// Trace: src/VX_cache_bank.sv:174:5
	assign req_idx_sel = (replay_valid ? replay_idx : core_req_idx);
	// Trace: src/VX_cache_bank.sv:175:5
	assign tag_sel = (init_valid | flush_valid ? (flush_valid ? flush_tag : {TAG_WIDTH {1'sb0}}) : (replay_valid ? replay_tag : (mem_rsp_valid ? mem_rsp_tag_s : core_req_tag)));
	// Trace: src/VX_cache_bank.sv:177:5
	assign flags_sel = (core_req_valid ? core_req_flags : {3 {1'sb0}});
	// Trace: src/VX_cache_bank.sv:178:5
	generate
		if (WRITE_ENABLE) begin : g_data_sel
			genvar _gv_i_195;
			for (_gv_i_195 = 0; _gv_i_195 < (8 * LINE_SIZE); _gv_i_195 = _gv_i_195 + 1) begin : g_i
				localparam i = _gv_i_195;
				if (i < (8 * WORD_SIZE)) begin : g_lo
					// Trace: src/VX_cache_bank.sv:181:17
					assign data_sel[i] = (replay_valid ? replay_data[i] : (mem_rsp_valid ? mem_rsp_data[i] : core_req_data[i]));
				end
				else begin : g_hi
					// Trace: src/VX_cache_bank.sv:183:17
					assign data_sel[i] = mem_rsp_data[i];
				end
			end
		end
		else begin : g_data_sel_ro
			// Trace: src/VX_cache_bank.sv:187:9
			assign data_sel = mem_rsp_data;
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:189:5
	generate
		if (1) begin : g_req_uuid_sel
			// Trace: src/VX_cache_bank.sv:190:9
			assign req_uuid_sel = tag_sel[TAG_WIDTH - 1-:VX_gpu_pkg_UUID_WIDTH];
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:194:5
	wire is_init_sel = init_valid;
	// Trace: src/VX_cache_bank.sv:195:5
	wire is_creq_sel = creq_enable || replay_enable;
	// Trace: src/VX_cache_bank.sv:196:5
	wire is_fill_sel = fill_enable;
	// Trace: src/VX_cache_bank.sv:197:5
	wire is_flush_sel = flush_enable;
	// Trace: src/VX_cache_bank.sv:198:5
	wire is_replay_sel = replay_enable;
	// Trace: src/VX_cache_bank.sv:199:5
	VX_pipe_register #(
		.DATAW(((((((((9 + ($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1)) + ((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS))) + (8 * LINE_SIZE)) + 1) + WORD_SIZE) + WORD_SEL_WIDTH) + REQ_SEL_WIDTH) + TAG_WIDTH) + MSHR_ADDR_WIDTH),
		.RESETW(1)
	) pipe_reg0(
		.clk(clk),
		.reset(reset),
		.enable(~pipe_stall),
		.data_in({valid_sel, is_init_sel, is_fill_sel, is_flush_sel, is_creq_sel, is_replay_sel, flags_sel, flush_way, addr_sel, data_sel, rw_sel, byteen_sel, word_idx_sel, req_idx_sel, tag_sel, replay_id}),
		.data_out({valid_st0, is_init_st0, is_fill_st0, is_flush_st0, is_creq_st0, is_replay_st0, flags_st0, flush_way_st0, addr_st0, data_st0, rw_st0, byteen_st0, word_idx_st0, req_idx_st0, tag_st0, replay_id_st0})
	);
	// Trace: src/VX_cache_bank.sv:209:5
	generate
		if (1) begin : g_req_uuid_st0
			// Trace: src/VX_cache_bank.sv:210:9
			assign req_uuid_st0 = tag_st0[TAG_WIDTH - 1-:VX_gpu_pkg_UUID_WIDTH];
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:214:5
	wire is_read_st0 = is_creq_st0 && ~rw_st0;
	// Trace: src/VX_cache_bank.sv:215:5
	wire is_write_st0 = is_creq_st0 && rw_st0;
	// Trace: src/VX_cache_bank.sv:216:5
	wire do_init_st0 = valid_st0 && is_init_st0;
	// Trace: src/VX_cache_bank.sv:217:5
	wire do_flush_st0 = valid_st0 && is_flush_st0;
	// Trace: src/VX_cache_bank.sv:218:5
	wire do_read_st0 = valid_st0 && is_read_st0;
	// Trace: src/VX_cache_bank.sv:219:5
	wire do_write_st0 = valid_st0 && is_write_st0;
	// Trace: src/VX_cache_bank.sv:220:5
	wire do_fill_st0 = valid_st0 && is_fill_st0;
	// Trace: src/VX_cache_bank.sv:221:5
	wire is_read_st1 = is_creq_st1 && ~rw_st1;
	// Trace: src/VX_cache_bank.sv:222:5
	wire is_write_st1 = is_creq_st1 && rw_st1;
	// Trace: src/VX_cache_bank.sv:223:5
	wire do_read_st1 = valid_st1 && is_read_st1;
	// Trace: src/VX_cache_bank.sv:224:5
	wire do_write_st1 = valid_st1 && is_write_st1;
	// Trace: src/VX_cache_bank.sv:225:5
	assign line_idx_sel = addr_sel[$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0];
	// Trace: src/VX_cache_bank.sv:226:5
	assign line_idx_st0 = addr_st0[$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0];
	// Trace: src/VX_cache_bank.sv:227:5
	assign line_tag_st0 = addr_st0[((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))];
	// Trace: src/VX_cache_bank.sv:228:5
	assign write_word_st0 = data_st0[(8 * WORD_SIZE) - 1:0];
	// Trace: src/VX_cache_bank.sv:229:5
	wire do_lookup_st0 = do_read_st0 || do_write_st0;
	// Trace: src/VX_cache_bank.sv:230:5
	wire do_lookup_st1 = do_read_st1 || do_write_st1;
	// Trace: src/VX_cache_bank.sv:231:5
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] victim_way_st0;
	// Trace: src/VX_cache_bank.sv:232:5
	wire [NUM_WAYS - 1:0] tag_matches_st0;
	// Trace: src/VX_cache_bank.sv:233:5
	VX_cache_repl #(
		.CACHE_SIZE(CACHE_SIZE),
		.LINE_SIZE(LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.NUM_WAYS(NUM_WAYS),
		.REPL_POLICY(REPL_POLICY)
	) cache_repl(
		.clk(clk),
		.reset(reset),
		.stall(pipe_stall),
		.init(do_init_st0),
		.lookup_valid(do_lookup_st1 && ~pipe_stall),
		.lookup_hit(is_hit_st1),
		.lookup_line(line_idx_st1),
		.lookup_way(way_idx_st1),
		.repl_valid(do_fill_st0 && ~pipe_stall),
		.repl_line(line_idx_st0),
		.repl_way(victim_way_st0)
	);
	// Trace: src/VX_cache_bank.sv:252:5
	assign evict_way_st0 = (is_fill_st0 ? victim_way_st0 : flush_way_st0);
	// Trace: src/VX_cache_bank.sv:253:5
	VX_cache_tags #(
		.CACHE_SIZE(CACHE_SIZE),
		.LINE_SIZE(LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.NUM_WAYS(NUM_WAYS),
		.WORD_SIZE(WORD_SIZE),
		.WRITEBACK(WRITEBACK)
	) cache_tags(
		.clk(clk),
		.reset(reset),
		.stall(pipe_stall),
		.init(do_init_st0),
		.flush(do_flush_st0 && ~pipe_stall),
		.fill(do_fill_st0 && ~pipe_stall),
		.read(do_read_st0 && ~pipe_stall),
		.write(do_write_st0 && ~pipe_stall),
		.line_idx(line_idx_st0),
		.line_idx_n(line_idx_sel),
		.line_tag(line_tag_st0),
		.evict_way(evict_way_st0),
		.tag_matches(tag_matches_st0),
		.evict_dirty(is_dirty_st0),
		.evict_tag(evict_tag_st0)
	);
	// Trace: src/VX_cache_bank.sv:277:5
	wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] hit_idx_st0;
	// Trace: src/VX_cache_bank.sv:278:5
	VX_onehot_encoder #(.N(NUM_WAYS)) way_idx_enc(
		.data_in(tag_matches_st0),
		.data_out(hit_idx_st0),
		.valid_out()
	);
	// Trace: src/VX_cache_bank.sv:285:5
	assign way_idx_st0 = (is_creq_st0 ? hit_idx_st0 : evict_way_st0);
	// Trace: src/VX_cache_bank.sv:286:5
	assign is_hit_st0 = |tag_matches_st0;
	// Trace: src/VX_cache_bank.sv:287:5
	wire [MSHR_ADDR_WIDTH - 1:0] mshr_alloc_id_st0;
	// Trace: src/VX_cache_bank.sv:288:5
	assign mshr_id_st0 = (is_replay_st0 ? replay_id_st0 : mshr_alloc_id_st0);
	// Trace: src/VX_cache_bank.sv:289:5
	VX_pipe_register #(
		.DATAW((((((((((((11 + ($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1)) + (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))) + (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) + (8 * LINE_SIZE)) + WORD_SIZE) + WORD_SEL_WIDTH) + REQ_SEL_WIDTH) + TAG_WIDTH) + MSHR_ADDR_WIDTH) + MSHR_ADDR_WIDTH) + 1),
		.RESETW(1)
	) pipe_reg1(
		.clk(clk),
		.reset(reset),
		.enable(~pipe_stall),
		.data_in({valid_st0, is_fill_st0, is_flush_st0, is_creq_st0, is_replay_st0, is_dirty_st0, is_hit_st0, rw_st0, flags_st0, way_idx_st0, evict_tag_st0, line_tag_st0, line_idx_st0, data_st0, byteen_st0, word_idx_st0, req_idx_st0, tag_st0, mshr_id_st0, mshr_previd_st0, mshr_pending_st0}),
		.data_out({valid_st1, is_fill_st1, is_flush_st1, is_creq_st1, is_replay_st1, is_dirty_st1, is_hit_st1, rw_st1, flags_st1, way_idx_st1, evict_tag_st1, line_tag_st1, line_idx_st1, data_st1, byteen_st1, word_idx_st1, req_idx_st1, tag_st1, mshr_id_st1, mshr_previd_st1, mshr_pending_st1})
	);
	// Trace: src/VX_cache_bank.sv:299:5
	generate
		if (1) begin : g_req_uuid_st1
			// Trace: src/VX_cache_bank.sv:300:9
			assign req_uuid_st1 = tag_st1[TAG_WIDTH - 1-:VX_gpu_pkg_UUID_WIDTH];
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:304:5
	assign addr_st1 = {line_tag_st1, line_idx_st1};
	// Trace: src/VX_cache_bank.sv:305:5
	assign write_word_st1 = data_st1[(8 * WORD_SIZE) - 1:0];
	// Trace: src/VX_cache_bank.sv:306:5
	wire [((LINE_SIZE / WORD_SIZE) * (8 * WORD_SIZE)) - 1:0] read_data_st1;
	// Trace: src/VX_cache_bank.sv:307:5
	wire [LINE_SIZE - 1:0] evict_byteen_st1;
	// Trace: src/VX_cache_bank.sv:308:5
	VX_cache_data #(
		.CACHE_SIZE(CACHE_SIZE),
		.LINE_SIZE(LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.NUM_WAYS(NUM_WAYS),
		.WORD_SIZE(WORD_SIZE),
		.WRITE_ENABLE(WRITE_ENABLE),
		.WRITEBACK(WRITEBACK),
		.DIRTY_BYTES(DIRTY_BYTES)
	) cache_data(
		.clk(clk),
		.reset(reset),
		.init(do_init_st0),
		.fill(do_fill_st0 && ~pipe_stall),
		.flush(do_flush_st0 && ~pipe_stall),
		.read(do_read_st0 && ~pipe_stall),
		.write(do_write_st0 && ~pipe_stall),
		.evict_way(evict_way_st0),
		.tag_matches(tag_matches_st0),
		.line_idx(line_idx_st0),
		.fill_data(data_st0),
		.write_word(write_word_st0),
		.word_idx(word_idx_st0),
		.write_byteen(byteen_st0),
		.way_idx_r(way_idx_st1),
		.read_data(read_data_st1),
		.evict_byteen(evict_byteen_st1)
	);
	// Trace: src/VX_cache_bank.sv:336:5
	wire mshr_allocate_st0 = (valid_st0 && is_creq_st0) && ~is_replay_st0;
	// Trace: src/VX_cache_bank.sv:337:5
	wire mshr_finalize_st1 = (valid_st1 && is_creq_st1) && ~is_replay_st1;
	// Trace: src/VX_cache_bank.sv:338:5
	wire mshr_release_st1;
	// Trace: src/VX_cache_bank.sv:339:5
	generate
		if (WRITEBACK) begin : g_mshr_release
			// Trace: src/VX_cache_bank.sv:340:9
			assign mshr_release_st1 = is_hit_st1;
		end
		else begin : g_mshr_release_ro
			// Trace: src/VX_cache_bank.sv:342:9
			assign mshr_release_st1 = is_hit_st1 || (rw_st1 && ~mshr_pending_st1);
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:344:5
	wire mshr_release_fire = (mshr_finalize_st1 && mshr_release_st1) && ~pipe_stall;
	// Trace: src/VX_cache_bank.sv:345:5
	wire [1:0] mshr_dequeue;
	// Trace: src/VX_cache_bank.sv:346:5
	VX_popcount #(
		.N(2),
		.MODEL(1)
	) __pop_count_ex482(
		.data_in({replay_fire, mshr_release_fire}),
		.data_out(mshr_dequeue)
	);
	// Trace: src/VX_cache_bank.sv:353:5
	VX_pending_size #(
		.SIZE(MSHR_SIZE),
		.DECRW(2)
	) mshr_pending_size(
		.clk(clk),
		.reset(reset),
		.incr(core_req_fire),
		.decr(mshr_dequeue),
		.empty(mshr_empty),
		.alm_empty(),
		.full(mshr_alm_full),
		.alm_full(),
		.size()
	);
	// Trace: src/VX_cache_bank.sv:367:5
	VX_cache_mshr #(
		.INSTANCE_ID(""),
		.BANK_ID(BANK_ID),
		.LINE_SIZE(LINE_SIZE),
		.NUM_BANKS(NUM_BANKS),
		.MSHR_SIZE(MSHR_SIZE),
		.WRITEBACK(WRITEBACK),
		.DATA_WIDTH((((WORD_SEL_WIDTH + WORD_SIZE) + (8 * WORD_SIZE)) + TAG_WIDTH) + REQ_SEL_WIDTH)
	) cache_mshr(
		.clk(clk),
		.reset(reset),
		.deq_req_uuid(req_uuid_sel),
		.alc_req_uuid(req_uuid_st0),
		.fin_req_uuid(req_uuid_st1),
		.fill_valid(mem_rsp_fire),
		.fill_id(mem_rsp_id),
		.fill_addr(mem_rsp_addr),
		.dequeue_valid(replay_valid),
		.dequeue_addr(replay_addr),
		.dequeue_rw(replay_rw),
		.dequeue_data({replay_wsel, replay_byteen, replay_data, replay_tag, replay_idx}),
		.dequeue_id(replay_id),
		.dequeue_ready(replay_ready),
		.allocate_valid(mshr_allocate_st0 && ~pipe_stall),
		.allocate_addr(addr_st0),
		.allocate_rw(rw_st0),
		.allocate_data({word_idx_st0, byteen_st0, write_word_st0, tag_st0, req_idx_st0}),
		.allocate_id(mshr_alloc_id_st0),
		.allocate_pending(mshr_pending_st0),
		.allocate_previd(mshr_previd_st0),
		.allocate_ready(),
		.finalize_valid(mshr_finalize_st1 && ~pipe_stall),
		.finalize_is_release(mshr_release_st1),
		.finalize_is_pending(mshr_pending_st1),
		.finalize_id(mshr_id_st1),
		.finalize_previd(mshr_previd_st1)
	);
	// Trace: src/VX_cache_bank.sv:404:5
	wire crsp_queue_valid;
	wire crsp_queue_ready;
	// Trace: src/VX_cache_bank.sv:405:5
	wire [(8 * WORD_SIZE) - 1:0] crsp_queue_data;
	// Trace: src/VX_cache_bank.sv:406:5
	wire [REQ_SEL_WIDTH - 1:0] crsp_queue_idx;
	// Trace: src/VX_cache_bank.sv:407:5
	wire [TAG_WIDTH - 1:0] crsp_queue_tag;
	// Trace: src/VX_cache_bank.sv:408:5
	assign crsp_queue_valid = do_read_st1 && is_hit_st1;
	// Trace: src/VX_cache_bank.sv:409:5
	assign crsp_queue_idx = req_idx_st1;
	// Trace: src/VX_cache_bank.sv:410:5
	assign crsp_queue_data = read_data_st1[word_idx_st1 * (8 * WORD_SIZE)+:8 * WORD_SIZE];
	// Trace: src/VX_cache_bank.sv:411:5
	assign crsp_queue_tag = tag_st1;
	// Trace: src/VX_cache_bank.sv:412:5
	VX_elastic_buffer #(
		.DATAW((TAG_WIDTH + (8 * WORD_SIZE)) + REQ_SEL_WIDTH),
		.SIZE(CRSQ_SIZE),
		.OUT_REG(CORE_OUT_REG)
	) core_rsp_queue(
		.clk(clk),
		.reset(reset),
		.valid_in(crsp_queue_valid),
		.ready_in(crsp_queue_ready),
		.data_in({crsp_queue_tag, crsp_queue_data, crsp_queue_idx}),
		.data_out({core_rsp_tag, core_rsp_data, core_rsp_idx}),
		.valid_out(core_rsp_valid),
		.ready_out(core_rsp_ready)
	);
	// Trace: src/VX_cache_bank.sv:426:5
	assign crsp_queue_stall = crsp_queue_valid && ~crsp_queue_ready;
	// Trace: src/VX_cache_bank.sv:427:5
	wire mreq_queue_push;
	wire mreq_queue_pop;
	// Trace: src/VX_cache_bank.sv:428:5
	wire [(8 * LINE_SIZE) - 1:0] mreq_queue_data;
	// Trace: src/VX_cache_bank.sv:429:5
	wire [LINE_SIZE - 1:0] mreq_queue_byteen;
	// Trace: src/VX_cache_bank.sv:430:5
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] mreq_queue_addr;
	// Trace: src/VX_cache_bank.sv:431:5
	wire [MEM_TAG_WIDTH - 1:0] mreq_queue_tag;
	// Trace: src/VX_cache_bank.sv:432:5
	wire mreq_queue_rw;
	// Trace: src/VX_cache_bank.sv:433:5
	wire [2:0] mreq_queue_flags;
	// Trace: src/VX_cache_bank.sv:434:5
	wire is_fill_or_flush_st1 = is_fill_st1 || (is_flush_st1 && WRITEBACK);
	// Trace: src/VX_cache_bank.sv:435:5
	wire do_fill_or_flush_st1 = valid_st1 && is_fill_or_flush_st1;
	// Trace: src/VX_cache_bank.sv:436:5
	wire do_writeback_st1 = do_fill_or_flush_st1 && is_dirty_st1;
	// Trace: src/VX_cache_bank.sv:437:5
	wire [((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS)) - 1:0] evict_addr_st1 = {evict_tag_st1, line_idx_st1};
	// Trace: src/VX_cache_bank.sv:438:5
	generate
		if (WRITE_ENABLE) begin : g_mreq_queue
			if (WRITEBACK) begin : g_wb
				if (DIRTY_BYTES) begin : g_dirty_bytes
					// Trace: src/VX_cache_bank.sv:441:17
					wire has_dirty_bytes = |evict_byteen_st1;
				end
				// Trace: src/VX_cache_bank.sv:443:13
				assign mreq_queue_push = (((do_lookup_st1 && ~is_hit_st1) && ~mshr_pending_st1) || do_writeback_st1) && ~pipe_stall;
				// Trace: src/VX_cache_bank.sv:446:13
				assign mreq_queue_addr = (is_fill_or_flush_st1 ? evict_addr_st1 : addr_st1);
				// Trace: src/VX_cache_bank.sv:447:13
				assign mreq_queue_rw = is_fill_or_flush_st1;
				// Trace: src/VX_cache_bank.sv:448:13
				assign mreq_queue_data = read_data_st1;
				// Trace: src/VX_cache_bank.sv:449:13
				assign mreq_queue_byteen = (is_fill_or_flush_st1 ? evict_byteen_st1 : {LINE_SIZE {1'sb1}});
			end
			else begin : g_wt
				// Trace: src/VX_cache_bank.sv:451:13
				wire [LINE_SIZE - 1:0] line_byteen;
				// Trace: src/VX_cache_bank.sv:452:13
				VX_demux #(
					.DATAW(WORD_SIZE),
					.N(LINE_SIZE / WORD_SIZE)
				) byteen_demux(
					.sel_in(word_idx_st1),
					.data_in(byteen_st1),
					.data_out(line_byteen)
				);
				// Trace: src/VX_cache_bank.sv:460:13
				assign mreq_queue_push = (((do_read_st1 && ~is_hit_st1) && ~mshr_pending_st1) || do_write_st1) && ~pipe_stall;
				// Trace: src/VX_cache_bank.sv:463:13
				assign mreq_queue_addr = addr_st1;
				// Trace: src/VX_cache_bank.sv:464:13
				assign mreq_queue_rw = rw_st1;
				// Trace: src/VX_cache_bank.sv:465:13
				assign mreq_queue_data = {LINE_SIZE / WORD_SIZE {write_word_st1}};
				// Trace: src/VX_cache_bank.sv:466:13
				assign mreq_queue_byteen = (rw_st1 ? line_byteen : {LINE_SIZE {1'sb1}});
			end
		end
		else begin : g_mreq_queue_ro
			// Trace: src/VX_cache_bank.sv:469:9
			assign mreq_queue_push = ((do_read_st1 && ~is_hit_st1) && ~mshr_pending_st1) && ~pipe_stall;
			// Trace: src/VX_cache_bank.sv:471:9
			assign mreq_queue_addr = addr_st1;
			// Trace: src/VX_cache_bank.sv:472:9
			assign mreq_queue_rw = 0;
			// Trace: src/VX_cache_bank.sv:473:9
			assign mreq_queue_data = 1'sb0;
			// Trace: src/VX_cache_bank.sv:474:9
			assign mreq_queue_byteen = 1'sb1;
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:476:5
	generate
		if (1) begin : g_mreq_queue_tag_uuid
			// Trace: src/VX_cache_bank.sv:477:9
			assign mreq_queue_tag = {req_uuid_st1, mshr_id_st1};
		end
	endgenerate
	// Trace: src/VX_cache_bank.sv:481:5
	assign mreq_queue_pop = mem_req_valid && mem_req_ready;
	// Trace: src/VX_cache_bank.sv:482:5
	assign mreq_queue_flags = flags_st1;
	// Trace: src/VX_cache_bank.sv:483:5
	VX_fifo_queue #(
		.DATAW(((((1 + ((32 - $clog2(LINE_SIZE)) - $clog2(NUM_BANKS))) + LINE_SIZE) + (8 * LINE_SIZE)) + MEM_TAG_WIDTH) + VX_gpu_pkg_MEM_FLAGS_WIDTH),
		.DEPTH(MREQ_SIZE),
		.ALM_FULL(MREQ_SIZE - PIPELINE_STAGES),
		.OUT_REG(MEM_OUT_REG)
	) mem_req_queue(
		.clk(clk),
		.reset(reset),
		.push(mreq_queue_push),
		.pop(mreq_queue_pop),
		.data_in({mreq_queue_rw, mreq_queue_addr, mreq_queue_byteen, mreq_queue_data, mreq_queue_tag, mreq_queue_flags}),
		.data_out({mem_req_rw, mem_req_addr, mem_req_byteen, mem_req_data, mem_req_tag, mem_req_flags}),
		.empty(mreq_queue_empty),
		.alm_full(mreq_queue_alm_full),
		.full(),
		.alm_empty(),
		.size()
	);
	// Trace: src/VX_cache_bank.sv:501:5
	assign mem_req_valid = ~mreq_queue_empty;
endmodule
// removed interface: VX_scoreboard_if
// removed module with interface ports: VX_local_mem
module VX_stream_switch (
	clk,
	reset,
	sel_in,
	valid_in,
	data_in,
	ready_in,
	valid_out,
	data_out,
	ready_out
);
	// Trace: src/VX_stream_switch.sv:2:15
	parameter NUM_INPUTS = 1;
	// Trace: src/VX_stream_switch.sv:3:15
	parameter NUM_OUTPUTS = 1;
	// Trace: src/VX_stream_switch.sv:4:15
	parameter DATAW = 1;
	// Trace: src/VX_stream_switch.sv:5:15
	parameter OUT_BUF = 0;
	// Trace: src/VX_stream_switch.sv:6:15
	parameter NUM_REQS = (NUM_INPUTS > NUM_OUTPUTS ? ((NUM_INPUTS + NUM_OUTPUTS) - 1) / NUM_OUTPUTS : ((NUM_OUTPUTS + NUM_INPUTS) - 1) / NUM_INPUTS);
	// Trace: src/VX_stream_switch.sv:7:15
	parameter SEL_COUNT = (NUM_INPUTS < NUM_OUTPUTS ? NUM_INPUTS : NUM_OUTPUTS);
	// Trace: src/VX_stream_switch.sv:8:15
	parameter LOG_NUM_REQS = $clog2(NUM_REQS);
	// Trace: src/VX_stream_switch.sv:10:5
	input wire clk;
	// Trace: src/VX_stream_switch.sv:11:5
	input wire reset;
	// Trace: src/VX_stream_switch.sv:12:5
	input wire [(SEL_COUNT * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)) - 1:0] sel_in;
	// Trace: src/VX_stream_switch.sv:13:5
	input wire [NUM_INPUTS - 1:0] valid_in;
	// Trace: src/VX_stream_switch.sv:14:5
	input wire [(NUM_INPUTS * DATAW) - 1:0] data_in;
	// Trace: src/VX_stream_switch.sv:15:5
	output wire [NUM_INPUTS - 1:0] ready_in;
	// Trace: src/VX_stream_switch.sv:16:5
	output wire [NUM_OUTPUTS - 1:0] valid_out;
	// Trace: src/VX_stream_switch.sv:17:5
	output wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out;
	// Trace: src/VX_stream_switch.sv:18:5
	input wire [NUM_OUTPUTS - 1:0] ready_out;
	// Trace: src/VX_stream_switch.sv:20:5
	wire [NUM_OUTPUTS - 1:0] valid_out_w;
	// Trace: src/VX_stream_switch.sv:21:5
	wire [(NUM_OUTPUTS * DATAW) - 1:0] data_out_w;
	// Trace: src/VX_stream_switch.sv:22:5
	wire [NUM_OUTPUTS - 1:0] ready_out_w;
	// Trace: src/VX_stream_switch.sv:23:5
	function automatic signed [LOG_NUM_REQS - 1:0] sv2v_cast_76B5F_signed;
		input reg signed [LOG_NUM_REQS - 1:0] inp;
		sv2v_cast_76B5F_signed = inp;
	endfunction
	generate
		if (NUM_INPUTS > NUM_OUTPUTS) begin : g_input_select
			genvar _gv_o_9;
			for (_gv_o_9 = 0; _gv_o_9 < NUM_OUTPUTS; _gv_o_9 = _gv_o_9 + 1) begin : g_out_buf
				localparam o = _gv_o_9;
				// Trace: src/VX_stream_switch.sv:25:13
				wire [NUM_REQS - 1:0] valid_in_w;
				// Trace: src/VX_stream_switch.sv:26:13
				wire [(NUM_REQS * DATAW) - 1:0] data_in_w;
				// Trace: src/VX_stream_switch.sv:27:13
				reg [NUM_REQS - 1:0] ready_in_w;
				genvar _gv_r_11;
				for (_gv_r_11 = 0; _gv_r_11 < NUM_REQS; _gv_r_11 = _gv_r_11 + 1) begin : g_r
					localparam r = _gv_r_11;
					// Trace: src/VX_stream_switch.sv:29:17
					localparam i = (r * NUM_OUTPUTS) + o;
					if (i < NUM_INPUTS) begin : g_valid
						// Trace: src/VX_stream_switch.sv:31:21
						assign valid_in_w[r] = valid_in[i];
						// Trace: src/VX_stream_switch.sv:32:21
						assign data_in_w[r * DATAW+:DATAW] = data_in[i * DATAW+:DATAW];
						// Trace: src/VX_stream_switch.sv:33:21
						assign ready_in[i] = ready_in_w[r];
					end
					else begin : g_padding
						// Trace: src/VX_stream_switch.sv:35:21
						assign valid_in_w[r] = 0;
						// Trace: src/VX_stream_switch.sv:36:21
						assign data_in_w[r * DATAW+:DATAW] = 1'sb0;
					end
				end
				// Trace: src/VX_stream_switch.sv:39:13
				assign valid_out_w[o] = valid_in_w[sel_in[o * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)+:(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)]];
				// Trace: src/VX_stream_switch.sv:40:13
				assign data_out_w[o * DATAW+:DATAW] = data_in_w[sel_in[o * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)+:(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)] * DATAW+:DATAW];
				// Trace: src/VX_stream_switch.sv:41:13
				always @(*) begin
					// Trace: src/VX_stream_switch.sv:42:17
					ready_in_w = 1'sb0;
					// Trace: src/VX_stream_switch.sv:43:17
					begin : sv2v_autoblock_1
						// Trace: src/VX_stream_switch.sv:43:22
						integer o;
						// Trace: src/VX_stream_switch.sv:43:22
						for (o = 0; o < NUM_OUTPUTS; o = o + 1)
							begin
								// Trace: src/VX_stream_switch.sv:44:21
								ready_in_w[sel_in[o * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)+:(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)]] = ready_out_w[o];
							end
					end
				end
			end
		end
		else if (NUM_OUTPUTS > NUM_INPUTS) begin : g_output_select
			genvar _gv_i_203;
			for (_gv_i_203 = 0; _gv_i_203 < NUM_INPUTS; _gv_i_203 = _gv_i_203 + 1) begin : g_out_buf
				localparam i = _gv_i_203;
				// Trace: src/VX_stream_switch.sv:50:13
				wire [NUM_REQS - 1:0] ready_out_s;
				genvar _gv_r_12;
				for (_gv_r_12 = 0; _gv_r_12 < NUM_REQS; _gv_r_12 = _gv_r_12 + 1) begin : g_r
					localparam r = _gv_r_12;
					// Trace: src/VX_stream_switch.sv:52:17
					localparam o = (r * NUM_INPUTS) + i;
					if (o < NUM_OUTPUTS) begin : g_valid
						// Trace: src/VX_stream_switch.sv:54:21
						assign valid_out_w[o] = valid_in[i] && (sel_in[i * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)+:(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)] == sv2v_cast_76B5F_signed(r));
						// Trace: src/VX_stream_switch.sv:55:21
						assign data_out_w[o * DATAW+:DATAW] = data_in[i * DATAW+:DATAW];
						// Trace: src/VX_stream_switch.sv:56:21
						assign ready_out_s[r] = ready_out_w[o];
					end
					else begin : g_padding
						// Trace: src/VX_stream_switch.sv:58:21
						assign ready_out_s[r] = 1'sb0;
					end
				end
				// Trace: src/VX_stream_switch.sv:61:13
				assign ready_in[i] = ready_out_s[sel_in[i * (LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)+:(LOG_NUM_REQS > 0 ? LOG_NUM_REQS : 1)]];
			end
		end
		else begin : g_passthru
			genvar _gv_i_204;
			for (_gv_i_204 = 0; _gv_i_204 < NUM_OUTPUTS; _gv_i_204 = _gv_i_204 + 1) begin : g_out_buf
				localparam i = _gv_i_204;
				// Trace: src/VX_stream_switch.sv:65:13
				assign valid_out_w[i] = valid_in[i];
				// Trace: src/VX_stream_switch.sv:66:13
				assign data_out_w[i * DATAW+:DATAW] = data_in[i * DATAW+:DATAW];
				// Trace: src/VX_stream_switch.sv:67:13
				assign ready_in[i] = ready_out_w[i];
			end
		end
	endgenerate
	// Trace: src/VX_stream_switch.sv:70:5
	genvar _gv_o_10;
	generate
		for (_gv_o_10 = 0; _gv_o_10 < NUM_OUTPUTS; _gv_o_10 = _gv_o_10 + 1) begin : g_out_buf
			localparam o = _gv_o_10;
			// Trace: src/VX_stream_switch.sv:71:9
			VX_elastic_buffer #(
				.DATAW(DATAW),
				.SIZE(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : 2)),
				.OUT_REG(((OUT_BUF & 7) < 2 ? OUT_BUF & 7 : (OUT_BUF & 7) - 2))
			) out_buf(
				.clk(clk),
				.reset(reset),
				.valid_in(valid_out_w[o]),
				.data_in(data_out_w[o * DATAW+:DATAW]),
				.ready_in(ready_out_w[o]),
				.valid_out(valid_out[o]),
				.data_out(data_out[o * DATAW+:DATAW]),
				.ready_out(ready_out[o])
			);
		end
	endgenerate
endmodule
module VX_pending_size (
	clk,
	reset,
	incr,
	decr,
	empty,
	alm_empty,
	full,
	alm_full,
	size
);
	// Trace: src/VX_pending_size.sv:2:15
	parameter SIZE = 1;
	// Trace: src/VX_pending_size.sv:3:15
	parameter INCRW = 1;
	// Trace: src/VX_pending_size.sv:4:15
	parameter DECRW = 1;
	// Trace: src/VX_pending_size.sv:5:15
	parameter ALM_FULL = SIZE - 1;
	// Trace: src/VX_pending_size.sv:6:15
	parameter ALM_EMPTY = 1;
	// Trace: src/VX_pending_size.sv:7:15
	parameter SIZEW = $clog2(SIZE + 1);
	// Trace: src/VX_pending_size.sv:9:5
	input wire clk;
	// Trace: src/VX_pending_size.sv:10:5
	input wire reset;
	// Trace: src/VX_pending_size.sv:11:5
	input wire [INCRW - 1:0] incr;
	// Trace: src/VX_pending_size.sv:12:5
	input wire [DECRW - 1:0] decr;
	// Trace: src/VX_pending_size.sv:13:5
	output wire empty;
	// Trace: src/VX_pending_size.sv:14:5
	output wire alm_empty;
	// Trace: src/VX_pending_size.sv:15:5
	output wire full;
	// Trace: src/VX_pending_size.sv:16:5
	output wire alm_full;
	// Trace: src/VX_pending_size.sv:17:5
	output wire [SIZEW - 1:0] size;
	// Trace: src/VX_pending_size.sv:19:5
	function automatic signed [SIZEW - 1:0] sv2v_cast_33A93_signed;
		input reg signed [SIZEW - 1:0] inp;
		sv2v_cast_33A93_signed = inp;
	endfunction
	generate
		if (SIZE == 1) begin : g_size_eq1
			// Trace: src/VX_pending_size.sv:20:9
			reg size_r;
			// Trace: src/VX_pending_size.sv:21:9
			always @(posedge clk)
				// Trace: src/VX_pending_size.sv:22:13
				if (reset)
					// Trace: src/VX_pending_size.sv:23:17
					size_r <= 1'sb0;
				else
					// Trace: src/VX_pending_size.sv:25:17
					if (incr) begin
						begin
							// Trace: src/VX_pending_size.sv:26:21
							if (~decr)
								// Trace: src/VX_pending_size.sv:27:25
								size_r <= 1;
						end
					end
					else if (decr)
						// Trace: src/VX_pending_size.sv:30:21
						size_r <= 1'sb0;
			// Trace: src/VX_pending_size.sv:34:9
			assign empty = size_r == 0;
			// Trace: src/VX_pending_size.sv:35:9
			assign full = size_r != 0;
			// Trace: src/VX_pending_size.sv:36:9
			assign alm_empty = 1'b1;
			// Trace: src/VX_pending_size.sv:37:9
			assign alm_full = 1'b1;
			// Trace: src/VX_pending_size.sv:38:9
			assign size = size_r;
		end
		else begin : g_size_gt1
			// Trace: src/VX_pending_size.sv:40:9
			reg empty_r;
			reg alm_empty_r;
			// Trace: src/VX_pending_size.sv:41:9
			reg full_r;
			reg alm_full_r;
			if ((INCRW != 1) || (DECRW != 1)) begin : g_wide_step
				// Trace: src/VX_pending_size.sv:43:13
				localparam DELTAW = (SIZEW < ((INCRW > DECRW ? INCRW : DECRW) + 1) ? SIZEW : (INCRW > DECRW ? INCRW : DECRW) + 1);
				// Trace: src/VX_pending_size.sv:44:13
				wire [SIZEW - 1:0] size_n;
				reg [SIZEW - 1:0] size_r;
				// Trace: src/VX_pending_size.sv:45:13
				function automatic [DELTAW - 1:0] sv2v_cast_B4011;
					input reg [DELTAW - 1:0] inp;
					sv2v_cast_B4011 = inp;
				endfunction
				wire [DELTAW - 1:0] delta = sv2v_cast_B4011(incr) - sv2v_cast_B4011(decr);
				// Trace: src/VX_pending_size.sv:46:13
				assign size_n = $signed(size_r) + sv2v_cast_33A93_signed($signed(delta));
				// Trace: src/VX_pending_size.sv:47:13
				always @(posedge clk)
					// Trace: src/VX_pending_size.sv:48:17
					if (reset) begin
						// Trace: src/VX_pending_size.sv:49:21
						empty_r <= 1;
						// Trace: src/VX_pending_size.sv:50:21
						full_r <= 0;
						// Trace: src/VX_pending_size.sv:51:21
						alm_empty_r <= 1;
						// Trace: src/VX_pending_size.sv:52:21
						alm_full_r <= 0;
						// Trace: src/VX_pending_size.sv:53:21
						size_r <= 1'sb0;
					end
					else begin
						// Trace: src/VX_pending_size.sv:55:21
						// Trace: src/VX_pending_size.sv:57:21
						empty_r <= size_n == sv2v_cast_33A93_signed(0);
						// Trace: src/VX_pending_size.sv:58:21
						full_r <= size_n == sv2v_cast_33A93_signed(SIZE);
						// Trace: src/VX_pending_size.sv:59:21
						alm_empty_r <= size_n <= sv2v_cast_33A93_signed(ALM_EMPTY);
						// Trace: src/VX_pending_size.sv:60:21
						alm_full_r <= size_n >= sv2v_cast_33A93_signed(ALM_FULL);
						// Trace: src/VX_pending_size.sv:61:21
						size_r <= size_n;
					end
				// Trace: src/VX_pending_size.sv:64:13
				assign size = size_r;
			end
			else begin : g_single_step
				// Trace: src/VX_pending_size.sv:66:13
				localparam ADDRW = (SIZE > 1 ? $clog2(SIZE) : 1);
				// Trace: src/VX_pending_size.sv:67:13
				reg [ADDRW - 1:0] used_r;
				// Trace: src/VX_pending_size.sv:68:13
				function automatic signed [ADDRW - 1:0] sv2v_cast_8BB5D_signed;
					input reg signed [ADDRW - 1:0] inp;
					sv2v_cast_8BB5D_signed = inp;
				endfunction
				wire is_alm_empty = used_r == sv2v_cast_8BB5D_signed(ALM_EMPTY);
				// Trace: src/VX_pending_size.sv:69:13
				wire is_alm_empty_n = used_r == sv2v_cast_8BB5D_signed(ALM_EMPTY + 1);
				// Trace: src/VX_pending_size.sv:70:13
				wire is_alm_full = used_r == sv2v_cast_8BB5D_signed(ALM_FULL);
				// Trace: src/VX_pending_size.sv:71:13
				wire is_alm_full_n = used_r == sv2v_cast_8BB5D_signed(ALM_FULL - 1);
				// Trace: src/VX_pending_size.sv:72:13
				always @(posedge clk)
					// Trace: src/VX_pending_size.sv:73:17
					if (reset) begin
						// Trace: src/VX_pending_size.sv:74:21
						alm_empty_r <= 1;
						// Trace: src/VX_pending_size.sv:75:21
						alm_full_r <= 0;
					end
					else
						// Trace: src/VX_pending_size.sv:77:21
						if (incr) begin
							begin
								// Trace: src/VX_pending_size.sv:78:25
								if (~decr) begin
									// Trace: src/VX_pending_size.sv:79:29
									if (is_alm_empty)
										// Trace: src/VX_pending_size.sv:80:33
										alm_empty_r <= 0;
									if (is_alm_full_n)
										// Trace: src/VX_pending_size.sv:82:33
										alm_full_r <= 1;
								end
							end
						end
						else if (decr) begin
							// Trace: src/VX_pending_size.sv:85:25
							if (is_alm_full)
								// Trace: src/VX_pending_size.sv:86:29
								alm_full_r <= 0;
							if (is_alm_empty_n)
								// Trace: src/VX_pending_size.sv:88:29
								alm_empty_r <= 1;
						end
				if (SIZE > 2) begin : g_size_gt2
					// Trace: src/VX_pending_size.sv:93:17
					function automatic signed [ADDRW - 1:0] sv2v_cast_8BB5D_signed;
						input reg signed [ADDRW - 1:0] inp;
						sv2v_cast_8BB5D_signed = inp;
					endfunction
					wire is_empty_n = used_r == sv2v_cast_8BB5D_signed(1);
					// Trace: src/VX_pending_size.sv:94:17
					wire is_full_n = used_r == sv2v_cast_8BB5D_signed(SIZE - 1);
					// Trace: src/VX_pending_size.sv:95:17
					wire [1:0] delta = {~incr & decr, incr ^ decr};
					// Trace: src/VX_pending_size.sv:96:17
					always @(posedge clk)
						// Trace: src/VX_pending_size.sv:97:21
						if (reset) begin
							// Trace: src/VX_pending_size.sv:98:25
							empty_r <= 1;
							// Trace: src/VX_pending_size.sv:99:25
							full_r <= 0;
							// Trace: src/VX_pending_size.sv:100:25
							used_r <= 1'sb0;
						end
						else begin
							// Trace: src/VX_pending_size.sv:102:25
							if (incr) begin
								begin
									// Trace: src/VX_pending_size.sv:103:29
									if (~decr) begin
										// Trace: src/VX_pending_size.sv:104:33
										empty_r <= 0;
										// Trace: src/VX_pending_size.sv:105:33
										if (is_full_n)
											// Trace: src/VX_pending_size.sv:106:37
											full_r <= 1;
									end
								end
							end
							else if (decr) begin
								// Trace: src/VX_pending_size.sv:109:29
								full_r <= 0;
								// Trace: src/VX_pending_size.sv:110:29
								if (is_empty_n)
									// Trace: src/VX_pending_size.sv:111:33
									empty_r <= 1;
							end
							// Trace: src/VX_pending_size.sv:113:25
							begin : sv2v_autoblock_1
								reg signed [ADDRW - 1:0] sv2v_tmp_cast;
								sv2v_tmp_cast = $signed(delta);
								used_r <= $signed(used_r) + sv2v_tmp_cast;
							end
						end
				end
				else begin : g_size_eq2
					// Trace: src/VX_pending_size.sv:117:17
					always @(posedge clk)
						// Trace: src/VX_pending_size.sv:118:21
						if (reset) begin
							// Trace: src/VX_pending_size.sv:119:25
							empty_r <= 1;
							// Trace: src/VX_pending_size.sv:120:25
							full_r <= 0;
							// Trace: src/VX_pending_size.sv:121:25
							used_r <= 1'sb0;
						end
						else begin
							// Trace: src/VX_pending_size.sv:123:25
							empty_r <= (empty_r & ~incr) | ((~full_r & decr) & ~incr);
							// Trace: src/VX_pending_size.sv:124:25
							full_r <= ((~empty_r & incr) & ~decr) | (full_r & ~(decr ^ incr));
							// Trace: src/VX_pending_size.sv:125:25
							used_r <= used_r ^ (incr ^ decr);
						end
				end
				if (SIZE > 1) begin : g_sizeN
					if (SIZEW > ADDRW) begin : g_not_log2
						// Trace: src/VX_pending_size.sv:131:21
						assign size = {full_r, used_r};
					end
					else begin : g_log2
						// Trace: src/VX_pending_size.sv:133:21
						assign size = used_r;
					end
				end
				else begin : g_size1
					// Trace: src/VX_pending_size.sv:136:17
					assign size = full_r;
				end
			end
			// Trace: src/VX_pending_size.sv:139:9
			assign empty = empty_r;
			// Trace: src/VX_pending_size.sv:140:9
			assign full = full_r;
			// Trace: src/VX_pending_size.sv:141:9
			assign alm_empty = alm_empty_r;
			// Trace: src/VX_pending_size.sv:142:9
			assign alm_full = alm_full_r;
		end
	endgenerate
endmodule
// removed interface: VX_fetch_if
// removed interface: VX_commit_if
// removed module with interface ports: VX_core
module VX_dp_ram (
	clk,
	reset,
	read,
	write,
	wren,
	waddr,
	wdata,
	raddr,
	rdata
);
	// Trace: src/VX_dp_ram.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_dp_ram.sv:3:15
	parameter SIZE = 1;
	// Trace: src/VX_dp_ram.sv:4:15
	parameter WRENW = 1;
	// Trace: src/VX_dp_ram.sv:5:15
	parameter OUT_REG = 0;
	// Trace: src/VX_dp_ram.sv:6:15
	parameter LUTRAM = 0;
	// Trace: src/VX_dp_ram.sv:7:15
	parameter RDW_MODE = "W";
	// Trace: src/VX_dp_ram.sv:8:15
	parameter RADDR_REG = 0;
	// Trace: src/VX_dp_ram.sv:9:15
	parameter RADDR_RESET = 0;
	// Trace: src/VX_dp_ram.sv:10:15
	parameter RDW_ASSERT = 0;
	// Trace: src/VX_dp_ram.sv:11:15
	parameter RESET_RAM = 0;
	// Trace: src/VX_dp_ram.sv:12:15
	parameter INIT_ENABLE = 0;
	// Trace: src/VX_dp_ram.sv:13:15
	parameter INIT_FILE = "";
	// Trace: src/VX_dp_ram.sv:14:15
	parameter [DATAW - 1:0] INIT_VALUE = 0;
	// Trace: src/VX_dp_ram.sv:15:15
	parameter ADDRW = (SIZE > 1 ? $clog2(SIZE) : 1);
	// Trace: src/VX_dp_ram.sv:17:5
	input wire clk;
	// Trace: src/VX_dp_ram.sv:18:5
	input wire reset;
	// Trace: src/VX_dp_ram.sv:19:5
	input wire read;
	// Trace: src/VX_dp_ram.sv:20:5
	input wire write;
	// Trace: src/VX_dp_ram.sv:21:5
	input wire [WRENW - 1:0] wren;
	// Trace: src/VX_dp_ram.sv:22:5
	input wire [ADDRW - 1:0] waddr;
	// Trace: src/VX_dp_ram.sv:23:5
	input wire [DATAW - 1:0] wdata;
	// Trace: src/VX_dp_ram.sv:24:5
	input wire [ADDRW - 1:0] raddr;
	// Trace: src/VX_dp_ram.sv:25:5
	output wire [DATAW - 1:0] rdata;
	// Trace: src/VX_dp_ram.sv:27:5
	localparam WSELW = DATAW / WRENW;
	// Trace: src/VX_dp_ram.sv:28:5
	localparam FORCE_BRAM = !LUTRAM && ((((SIZE >= 64) || (DATAW >= 16)) || ((SIZE * DATAW) >= 512)) && ((SIZE * DATAW) >= 64));
	// Trace: src/VX_dp_ram.sv:29:5
	generate
		if (OUT_REG) begin : g_sync
			if (FORCE_BRAM) begin : g_bram
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:33:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:36:13
								initial begin
									// Trace: src/VX_dp_ram.sv:36:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:38:13
								initial begin
									// Trace: src/VX_dp_ram.sv:39:17
									begin : sv2v_autoblock_1
										// Trace: src/VX_dp_ram.sv:39:22
										integer i;
										// Trace: src/VX_dp_ram.sv:39:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:40:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:45:21
						reg [ADDRW - 1:0] raddr_r;
						// Trace: src/VX_dp_ram.sv:46:21
						always @(posedge clk) begin
							// Trace: src/VX_dp_ram.sv:47:29
							if (write)
								// Trace: src/VX_dp_ram.sv:48:33
								begin : sv2v_autoblock_2
									// Trace: src/VX_dp_ram.sv:48:38
									integer i;
									// Trace: src/VX_dp_ram.sv:48:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:49:37
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:50:41
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							if (read)
								// Trace: src/VX_dp_ram.sv:55:29
								raddr_r <= raddr;
						end
						// Trace: src/VX_dp_ram.sv:58:21
						assign rdata = ram[raddr_r];
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:60:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:63:13
								initial begin
									// Trace: src/VX_dp_ram.sv:63:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:65:13
								initial begin
									// Trace: src/VX_dp_ram.sv:66:17
									begin : sv2v_autoblock_3
										// Trace: src/VX_dp_ram.sv:66:22
										integer i;
										// Trace: src/VX_dp_ram.sv:66:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:67:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:72:21
						reg [ADDRW - 1:0] raddr_r;
						// Trace: src/VX_dp_ram.sv:73:21
						always @(posedge clk) begin
							// Trace: src/VX_dp_ram.sv:74:25
							if (write)
								// Trace: src/VX_dp_ram.sv:75:29
								ram[waddr] <= wdata;
							if (read)
								// Trace: src/VX_dp_ram.sv:78:29
								raddr_r <= raddr;
						end
						// Trace: src/VX_dp_ram.sv:81:21
						assign rdata = ram[raddr_r];
					end
				end
				else if (RDW_MODE == "R") begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:85:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:88:13
								initial begin
									// Trace: src/VX_dp_ram.sv:88:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:90:13
								initial begin
									// Trace: src/VX_dp_ram.sv:91:17
									begin : sv2v_autoblock_4
										// Trace: src/VX_dp_ram.sv:91:22
										integer i;
										// Trace: src/VX_dp_ram.sv:91:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:92:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:97:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_dp_ram.sv:98:21
						always @(posedge clk) begin
							// Trace: src/VX_dp_ram.sv:99:29
							if (write)
								// Trace: src/VX_dp_ram.sv:100:33
								begin : sv2v_autoblock_5
									// Trace: src/VX_dp_ram.sv:100:38
									integer i;
									// Trace: src/VX_dp_ram.sv:100:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:101:37
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:102:41
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							if (read)
								// Trace: src/VX_dp_ram.sv:107:29
								rdata_r <= ram[raddr];
						end
						// Trace: src/VX_dp_ram.sv:110:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:112:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:115:13
								initial begin
									// Trace: src/VX_dp_ram.sv:115:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:117:13
								initial begin
									// Trace: src/VX_dp_ram.sv:118:17
									begin : sv2v_autoblock_6
										// Trace: src/VX_dp_ram.sv:118:22
										integer i;
										// Trace: src/VX_dp_ram.sv:118:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:119:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:124:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_dp_ram.sv:125:21
						always @(posedge clk) begin
							// Trace: src/VX_dp_ram.sv:126:25
							if (write)
								// Trace: src/VX_dp_ram.sv:127:29
								ram[waddr] <= wdata;
							if (read)
								// Trace: src/VX_dp_ram.sv:130:29
								rdata_r <= ram[raddr];
						end
						// Trace: src/VX_dp_ram.sv:133:21
						assign rdata = rdata_r;
					end
				end
			end
			else begin : g_auto
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:139:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:142:13
								initial begin
									// Trace: src/VX_dp_ram.sv:142:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:144:13
								initial begin
									// Trace: src/VX_dp_ram.sv:145:17
									begin : sv2v_autoblock_7
										// Trace: src/VX_dp_ram.sv:145:22
										integer i;
										// Trace: src/VX_dp_ram.sv:145:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:146:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:151:21
						reg [ADDRW - 1:0] raddr_r;
						// Trace: src/VX_dp_ram.sv:152:21
						always @(posedge clk) begin
							// Trace: src/VX_dp_ram.sv:153:29
							if (write)
								// Trace: src/VX_dp_ram.sv:154:33
								begin : sv2v_autoblock_8
									// Trace: src/VX_dp_ram.sv:154:38
									integer i;
									// Trace: src/VX_dp_ram.sv:154:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:155:37
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:156:41
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							if (read)
								// Trace: src/VX_dp_ram.sv:161:29
								raddr_r <= raddr;
						end
						// Trace: src/VX_dp_ram.sv:164:21
						assign rdata = ram[raddr_r];
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:166:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:169:13
								initial begin
									// Trace: src/VX_dp_ram.sv:169:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:171:13
								initial begin
									// Trace: src/VX_dp_ram.sv:172:17
									begin : sv2v_autoblock_9
										// Trace: src/VX_dp_ram.sv:172:22
										integer i;
										// Trace: src/VX_dp_ram.sv:172:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:173:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:178:21
						reg [ADDRW - 1:0] raddr_r;
						// Trace: src/VX_dp_ram.sv:179:21
						always @(posedge clk) begin
							// Trace: src/VX_dp_ram.sv:180:25
							if (write)
								// Trace: src/VX_dp_ram.sv:181:29
								ram[waddr] <= wdata;
							if (read)
								// Trace: src/VX_dp_ram.sv:184:29
								raddr_r <= raddr;
						end
						// Trace: src/VX_dp_ram.sv:187:21
						assign rdata = ram[raddr_r];
					end
				end
				else if (RDW_MODE == "R") begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:191:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:194:13
								initial begin
									// Trace: src/VX_dp_ram.sv:194:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:196:13
								initial begin
									// Trace: src/VX_dp_ram.sv:197:17
									begin : sv2v_autoblock_10
										// Trace: src/VX_dp_ram.sv:197:22
										integer i;
										// Trace: src/VX_dp_ram.sv:197:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:198:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:203:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_dp_ram.sv:204:21
						always @(posedge clk) begin
							// Trace: src/VX_dp_ram.sv:205:29
							if (write)
								// Trace: src/VX_dp_ram.sv:206:33
								begin : sv2v_autoblock_11
									// Trace: src/VX_dp_ram.sv:206:38
									integer i;
									// Trace: src/VX_dp_ram.sv:206:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:207:37
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:208:41
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
							if (read)
								// Trace: src/VX_dp_ram.sv:213:29
								rdata_r <= ram[raddr];
						end
						// Trace: src/VX_dp_ram.sv:216:21
						assign rdata = rdata_r;
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:218:21
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:221:13
								initial begin
									// Trace: src/VX_dp_ram.sv:221:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:223:13
								initial begin
									// Trace: src/VX_dp_ram.sv:224:17
									begin : sv2v_autoblock_12
										// Trace: src/VX_dp_ram.sv:224:22
										integer i;
										// Trace: src/VX_dp_ram.sv:224:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:225:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:230:21
						reg [DATAW - 1:0] rdata_r;
						// Trace: src/VX_dp_ram.sv:231:21
						always @(posedge clk) begin
							// Trace: src/VX_dp_ram.sv:232:25
							if (write)
								// Trace: src/VX_dp_ram.sv:233:29
								ram[waddr] <= wdata;
							if (read)
								// Trace: src/VX_dp_ram.sv:236:29
								rdata_r <= ram[raddr];
						end
						// Trace: src/VX_dp_ram.sv:239:21
						assign rdata = rdata_r;
					end
				end
			end
		end
		else begin : g_async
			if (FORCE_BRAM) begin : g_bram
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:247:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:250:13
								initial begin
									// Trace: src/VX_dp_ram.sv:250:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:252:13
								initial begin
									// Trace: src/VX_dp_ram.sv:253:17
									begin : sv2v_autoblock_13
										// Trace: src/VX_dp_ram.sv:253:22
										integer i;
										// Trace: src/VX_dp_ram.sv:253:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:254:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:259:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:260:29
							if (write)
								// Trace: src/VX_dp_ram.sv:261:33
								begin : sv2v_autoblock_14
									// Trace: src/VX_dp_ram.sv:261:38
									integer i;
									// Trace: src/VX_dp_ram.sv:261:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:262:37
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:263:41
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_dp_ram.sv:268:21
						assign rdata = ram[raddr];
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:270:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:273:13
								initial begin
									// Trace: src/VX_dp_ram.sv:273:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:275:13
								initial begin
									// Trace: src/VX_dp_ram.sv:276:17
									begin : sv2v_autoblock_15
										// Trace: src/VX_dp_ram.sv:276:22
										integer i;
										// Trace: src/VX_dp_ram.sv:276:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:277:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:282:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:283:25
							if (write)
								// Trace: src/VX_dp_ram.sv:284:29
								ram[waddr] <= wdata;
						// Trace: src/VX_dp_ram.sv:287:21
						assign rdata = ram[raddr];
					end
				end
				else begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:291:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:294:13
								initial begin
									// Trace: src/VX_dp_ram.sv:294:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:296:13
								initial begin
									// Trace: src/VX_dp_ram.sv:297:17
									begin : sv2v_autoblock_16
										// Trace: src/VX_dp_ram.sv:297:22
										integer i;
										// Trace: src/VX_dp_ram.sv:297:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:298:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:303:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:304:29
							if (write)
								// Trace: src/VX_dp_ram.sv:305:33
								begin : sv2v_autoblock_17
									// Trace: src/VX_dp_ram.sv:305:38
									integer i;
									// Trace: src/VX_dp_ram.sv:305:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:306:37
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:307:41
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_dp_ram.sv:312:21
						assign rdata = ram[raddr];
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:314:23
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:317:13
								initial begin
									// Trace: src/VX_dp_ram.sv:317:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:319:13
								initial begin
									// Trace: src/VX_dp_ram.sv:320:17
									begin : sv2v_autoblock_18
										// Trace: src/VX_dp_ram.sv:320:22
										integer i;
										// Trace: src/VX_dp_ram.sv:320:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:321:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:326:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:327:25
							if (write)
								// Trace: src/VX_dp_ram.sv:328:29
								ram[waddr] <= wdata;
						// Trace: src/VX_dp_ram.sv:331:21
						assign rdata = ram[raddr];
					end
				end
			end
			else begin : g_auto
				if (RDW_MODE == "W") begin : g_write_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:337:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:340:13
								initial begin
									// Trace: src/VX_dp_ram.sv:340:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:342:13
								initial begin
									// Trace: src/VX_dp_ram.sv:343:17
									begin : sv2v_autoblock_19
										// Trace: src/VX_dp_ram.sv:343:22
										integer i;
										// Trace: src/VX_dp_ram.sv:343:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:344:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:349:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:350:29
							if (write)
								// Trace: src/VX_dp_ram.sv:351:33
								begin : sv2v_autoblock_20
									// Trace: src/VX_dp_ram.sv:351:38
									integer i;
									// Trace: src/VX_dp_ram.sv:351:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:352:37
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:353:41
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_dp_ram.sv:358:21
						assign rdata = ram[raddr];
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:360:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:363:13
								initial begin
									// Trace: src/VX_dp_ram.sv:363:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:365:13
								initial begin
									// Trace: src/VX_dp_ram.sv:366:17
									begin : sv2v_autoblock_21
										// Trace: src/VX_dp_ram.sv:366:22
										integer i;
										// Trace: src/VX_dp_ram.sv:366:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:367:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:372:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:373:25
							if (write)
								// Trace: src/VX_dp_ram.sv:374:29
								ram[waddr] <= wdata;
						// Trace: src/VX_dp_ram.sv:377:21
						assign rdata = ram[raddr];
					end
				end
				else begin : g_read_first
					if (WRENW != 1) begin : g_wren
						// Trace: src/VX_dp_ram.sv:381:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:384:13
								initial begin
									// Trace: src/VX_dp_ram.sv:384:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:386:13
								initial begin
									// Trace: src/VX_dp_ram.sv:387:17
									begin : sv2v_autoblock_22
										// Trace: src/VX_dp_ram.sv:387:22
										integer i;
										// Trace: src/VX_dp_ram.sv:387:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:388:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:393:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:394:29
							if (write)
								// Trace: src/VX_dp_ram.sv:395:33
								begin : sv2v_autoblock_23
									// Trace: src/VX_dp_ram.sv:395:38
									integer i;
									// Trace: src/VX_dp_ram.sv:395:38
									for (i = 0; i < WRENW; i = i + 1)
										begin
											// Trace: src/VX_dp_ram.sv:396:37
											if (wren[i])
												// Trace: src/VX_dp_ram.sv:397:41
												ram[waddr][i * WSELW+:WSELW] <= wdata[i * WSELW+:WSELW];
										end
								end
						// Trace: src/VX_dp_ram.sv:402:21
						assign rdata = ram[raddr];
					end
					else begin : g_no_wren
						// Trace: src/VX_dp_ram.sv:404:22
						reg [DATAW - 1:0] ram [0:SIZE - 1];
						if (INIT_ENABLE != 0) begin : g_init
							if (INIT_FILE != "") begin : g_file
								// Trace: src/VX_dp_ram.sv:407:13
								initial begin
									// Trace: src/VX_dp_ram.sv:407:21
									$readmemh(INIT_FILE, ram);
								end
							end
							else begin : g_value
								// Trace: src/VX_dp_ram.sv:409:13
								initial begin
									// Trace: src/VX_dp_ram.sv:410:17
									begin : sv2v_autoblock_24
										// Trace: src/VX_dp_ram.sv:410:22
										integer i;
										// Trace: src/VX_dp_ram.sv:410:22
										for (i = 0; i < SIZE; i = i + 1)
											begin : g_i
												// Trace: src/VX_dp_ram.sv:411:21
												ram[i] = INIT_VALUE;
											end
									end
								end
							end
						end
						// Trace: src/VX_dp_ram.sv:416:21
						always @(posedge clk)
							// Trace: src/VX_dp_ram.sv:417:25
							if (write)
								// Trace: src/VX_dp_ram.sv:418:29
								ram[waddr] <= wdata;
						// Trace: src/VX_dp_ram.sv:421:21
						assign rdata = ram[raddr];
					end
				end
			end
		end
	endgenerate
endmodule
// removed module with interface ports: VX_fetch
// removed module with interface ports: VX_operands
module VX_cache_tags (
	clk,
	reset,
	stall,
	init,
	flush,
	fill,
	read,
	write,
	line_idx,
	line_idx_n,
	line_tag,
	evict_way,
	tag_matches,
	evict_dirty,
	evict_tag
);
	// removed import VX_gpu_pkg::*;
	// Trace: src/VX_cache_tags.sv:2:15
	parameter CACHE_SIZE = 1024;
	// Trace: src/VX_cache_tags.sv:3:15
	parameter LINE_SIZE = 16;
	// Trace: src/VX_cache_tags.sv:4:15
	parameter NUM_BANKS = 1;
	// Trace: src/VX_cache_tags.sv:5:15
	parameter NUM_WAYS = 1;
	// Trace: src/VX_cache_tags.sv:6:15
	parameter WORD_SIZE = 1;
	// Trace: src/VX_cache_tags.sv:7:15
	parameter WRITEBACK = 0;
	// Trace: src/VX_cache_tags.sv:9:5
	input wire clk;
	// Trace: src/VX_cache_tags.sv:10:5
	input wire reset;
	// Trace: src/VX_cache_tags.sv:11:5
	input wire stall;
	// Trace: src/VX_cache_tags.sv:12:5
	input wire init;
	// Trace: src/VX_cache_tags.sv:13:5
	input wire flush;
	// Trace: src/VX_cache_tags.sv:14:5
	input wire fill;
	// Trace: src/VX_cache_tags.sv:15:5
	input wire read;
	// Trace: src/VX_cache_tags.sv:16:5
	input wire write;
	// Trace: src/VX_cache_tags.sv:17:5
	input wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] line_idx;
	// Trace: src/VX_cache_tags.sv:18:5
	input wire [$clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)) - 1:0] line_idx_n;
	// Trace: src/VX_cache_tags.sv:19:5
	input wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) - 1:0] line_tag;
	// Trace: src/VX_cache_tags.sv:20:5
	input wire [($clog2(NUM_WAYS) > 0 ? $clog2(NUM_WAYS) : 1) - 1:0] evict_way;
	// Trace: src/VX_cache_tags.sv:21:5
	output wire [NUM_WAYS - 1:0] tag_matches;
	// Trace: src/VX_cache_tags.sv:22:5
	output wire evict_dirty;
	// Trace: src/VX_cache_tags.sv:23:5
	output wire [(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) - 1:0] evict_tag;
	// Trace: src/VX_cache_tags.sv:25:5
	localparam TAG_WIDTH = (1 + WRITEBACK) + (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1));
	// Trace: src/VX_cache_tags.sv:26:5
	wire [(NUM_WAYS * (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))) - 1:0] read_tag;
	// Trace: src/VX_cache_tags.sv:27:5
	wire [NUM_WAYS - 1:0] read_valid;
	// Trace: src/VX_cache_tags.sv:28:5
	wire [NUM_WAYS - 1:0] read_dirty;
	// Trace: src/VX_cache_tags.sv:29:5
	generate
		if (WRITEBACK) begin : g_evict_tag_wb
			// Trace: src/VX_cache_tags.sv:30:9
			assign evict_dirty = read_dirty[evict_way];
			// Trace: src/VX_cache_tags.sv:31:9
			assign evict_tag = read_tag[evict_way * (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))+:((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)];
		end
		else begin : g_evict_tag_wt
			// Trace: src/VX_cache_tags.sv:33:9
			assign evict_dirty = 1'b0;
			// Trace: src/VX_cache_tags.sv:34:9
			assign evict_tag = 1'sb0;
		end
	endgenerate
	// Trace: src/VX_cache_tags.sv:36:5
	genvar _gv_i_208;
	generate
		for (_gv_i_208 = 0; _gv_i_208 < NUM_WAYS; _gv_i_208 = _gv_i_208 + 1) begin : g_tag_store
			localparam i = _gv_i_208;
			// Trace: src/VX_cache_tags.sv:37:9
			wire way_en = (NUM_WAYS == 1) || (evict_way == i);
			// Trace: src/VX_cache_tags.sv:38:9
			wire do_init = init;
			// Trace: src/VX_cache_tags.sv:39:9
			wire do_fill = fill && way_en;
			// Trace: src/VX_cache_tags.sv:40:9
			wire do_flush = flush && (!WRITEBACK || way_en);
			// Trace: src/VX_cache_tags.sv:41:9
			wire do_write = (WRITEBACK && write) && tag_matches[i];
			// Trace: src/VX_cache_tags.sv:42:9
			wire line_write = ((do_init || do_fill) || do_flush) || do_write;
			// Trace: src/VX_cache_tags.sv:43:9
			wire line_valid = fill || write;
			// Trace: src/VX_cache_tags.sv:44:9
			wire [TAG_WIDTH - 1:0] line_wdata;
			wire [TAG_WIDTH - 1:0] line_rdata;
			// Trace: src/VX_cache_tags.sv:45:9
			wire rdw_fill;
			wire rdw_write;
			// Trace: src/VX_cache_tags.sv:46:5
			VX_pipe_register #(
				.DATAW(1),
				.RESETW(1),
				.DEPTH(1)
			) __buffer_ex84(
				.clk(clk),
				.reset(reset),
				.enable(1'b1),
				.data_in(do_fill),
				.data_out(rdw_fill)
			);
			// Trace: src/VX_cache_tags.sv:57:5
			VX_pipe_register #(
				.DATAW(1),
				.RESETW(1),
				.DEPTH(1)
			) __buffer_ex85(
				.clk(clk),
				.reset(reset),
				.enable(1'b1),
				.data_in(do_write && (line_idx == line_idx_n)),
				.data_out(rdw_write)
			);
			if (WRITEBACK) begin : g_wdata
				// Trace: src/VX_cache_tags.sv:69:13
				assign line_wdata = {line_valid, write, line_tag};
				// Trace: src/VX_cache_tags.sv:70:13
				assign read_tag[i * (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))+:((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)] = line_rdata[0+:((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)];
				// Trace: src/VX_cache_tags.sv:71:13
				assign read_dirty[i] = line_rdata[((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)] || rdw_write;
				// Trace: src/VX_cache_tags.sv:72:13
				assign read_valid[i] = line_rdata[(((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)) + 1];
			end
			else begin : g_wdata
				// Trace: src/VX_cache_tags.sv:74:13
				assign line_wdata = {line_valid, line_tag};
				// Trace: src/VX_cache_tags.sv:75:13
				assign {read_valid[i], read_tag[i * (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))+:((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)]} = line_rdata;
				// Trace: src/VX_cache_tags.sv:76:13
				assign read_dirty[i] = 1'b0;
			end
			// Trace: src/VX_cache_tags.sv:78:9
			VX_dp_ram #(
				.DATAW(TAG_WIDTH),
				.SIZE((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS)),
				.OUT_REG(1),
				.RDW_MODE("R")
			) tag_store(
				.clk(clk),
				.reset(reset),
				.read(~stall),
				.write(line_write),
				.wren(1'b1),
				.waddr(line_idx),
				.raddr(line_idx_n),
				.wdata(line_wdata),
				.rdata(line_rdata)
			);
			// Trace: src/VX_cache_tags.sv:94:9
			assign tag_matches[i] = (read_valid[i] && (line_tag == read_tag[i * (((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1))+:((32 - $clog2(WORD_SIZE)) - 1) - ((((((0 + $clog2(LINE_SIZE / WORD_SIZE)) + 0) + $clog2(NUM_BANKS)) + 0) + $clog2((CACHE_SIZE / NUM_BANKS) / (LINE_SIZE * NUM_WAYS))) - 1)])) || rdw_fill;
		end
	endgenerate
endmodule
module VX_priority_arbiter (
	clk,
	reset,
	requests,
	grant_index,
	grant_onehot,
	grant_valid,
	grant_ready
);
	// Trace: src/VX_priority_arbiter.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_priority_arbiter.sv:3:15
	parameter STICKY = 0;
	// Trace: src/VX_priority_arbiter.sv:4:15
	parameter LOG_NUM_REQS = (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1);
	// Trace: src/VX_priority_arbiter.sv:6:5
	input wire clk;
	// Trace: src/VX_priority_arbiter.sv:7:5
	input wire reset;
	// Trace: src/VX_priority_arbiter.sv:8:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: src/VX_priority_arbiter.sv:9:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: src/VX_priority_arbiter.sv:10:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: src/VX_priority_arbiter.sv:11:5
	output wire grant_valid;
	// Trace: src/VX_priority_arbiter.sv:12:5
	input wire grant_ready;
	// Trace: src/VX_priority_arbiter.sv:14:5
	generate
		if (NUM_REQS == 1) begin : g_passthru
			// Trace: src/VX_priority_arbiter.sv:15:9
			assign grant_index = 1'sb0;
			// Trace: src/VX_priority_arbiter.sv:16:9
			assign grant_onehot = requests;
			// Trace: src/VX_priority_arbiter.sv:17:9
			assign grant_valid = requests[0];
		end
		else begin : g_encoder
			// Trace: src/VX_priority_arbiter.sv:19:9
			reg [NUM_REQS - 1:0] prev_grant;
			// Trace: src/VX_priority_arbiter.sv:20:9
			always @(posedge clk)
				// Trace: src/VX_priority_arbiter.sv:21:13
				if (reset)
					// Trace: src/VX_priority_arbiter.sv:22:17
					prev_grant <= 1'sb0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_priority_arbiter.sv:24:17
					prev_grant <= grant_onehot;
			// Trace: src/VX_priority_arbiter.sv:27:9
			wire retain_grant = (STICKY != 0) && |(prev_grant & requests);
			// Trace: src/VX_priority_arbiter.sv:28:9
			wire [NUM_REQS - 1:0] requests_w = (retain_grant ? prev_grant : requests);
			// Trace: src/VX_priority_arbiter.sv:29:9
			wire grant_valid_w;
			// Trace: src/VX_priority_arbiter.sv:30:9
			VX_priority_encoder #(.N(NUM_REQS)) grant_sel(
				.data_in(requests_w),
				.index_out(grant_index),
				.onehot_out(grant_onehot),
				.valid_out(grant_valid_w)
			);
			// Trace: src/VX_priority_arbiter.sv:38:9
			assign grant_valid = (STICKY != 0 ? |requests : grant_valid_w);
		end
	endgenerate
endmodule
module VX_cyclic_arbiter (
	clk,
	reset,
	requests,
	grant_index,
	grant_onehot,
	grant_valid,
	grant_ready
);
	// Trace: src/VX_cyclic_arbiter.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_cyclic_arbiter.sv:3:15
	parameter STICKY = 0;
	// Trace: src/VX_cyclic_arbiter.sv:4:15
	parameter LOG_NUM_REQS = (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1);
	// Trace: src/VX_cyclic_arbiter.sv:6:5
	input wire clk;
	// Trace: src/VX_cyclic_arbiter.sv:7:5
	input wire reset;
	// Trace: src/VX_cyclic_arbiter.sv:8:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: src/VX_cyclic_arbiter.sv:9:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: src/VX_cyclic_arbiter.sv:10:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: src/VX_cyclic_arbiter.sv:11:5
	output wire grant_valid;
	// Trace: src/VX_cyclic_arbiter.sv:12:5
	input wire grant_ready;
	// Trace: src/VX_cyclic_arbiter.sv:14:5
	function automatic signed [LOG_NUM_REQS - 1:0] sv2v_cast_76B5F_signed;
		input reg signed [LOG_NUM_REQS - 1:0] inp;
		sv2v_cast_76B5F_signed = inp;
	endfunction
	generate
		if (NUM_REQS == 1) begin : g_passthru
			// Trace: src/VX_cyclic_arbiter.sv:15:9
			assign grant_index = 1'sb0;
			// Trace: src/VX_cyclic_arbiter.sv:16:9
			assign grant_onehot = requests;
			// Trace: src/VX_cyclic_arbiter.sv:17:9
			assign grant_valid = requests[0];
		end
		else begin : g_arbiter
			// Trace: src/VX_cyclic_arbiter.sv:19:9
			localparam IS_POW2 = (1 << LOG_NUM_REQS) == NUM_REQS;
			// Trace: src/VX_cyclic_arbiter.sv:20:9
			wire [LOG_NUM_REQS - 1:0] grant_index_um;
			// Trace: src/VX_cyclic_arbiter.sv:21:9
			wire [NUM_REQS - 1:0] grant_onehot_w;
			wire [NUM_REQS - 1:0] grant_onehot_um;
			// Trace: src/VX_cyclic_arbiter.sv:22:9
			reg [LOG_NUM_REQS - 1:0] grant_index_r;
			// Trace: src/VX_cyclic_arbiter.sv:23:9
			reg [NUM_REQS - 1:0] prev_grant;
			// Trace: src/VX_cyclic_arbiter.sv:24:9
			always @(posedge clk)
				// Trace: src/VX_cyclic_arbiter.sv:25:13
				if (reset)
					// Trace: src/VX_cyclic_arbiter.sv:26:17
					prev_grant <= 1'sb0;
				else if (grant_valid && grant_ready)
					// Trace: src/VX_cyclic_arbiter.sv:28:17
					prev_grant <= grant_onehot;
			// Trace: src/VX_cyclic_arbiter.sv:31:9
			wire retain_grant = (STICKY != 0) && |(prev_grant & requests);
			// Trace: src/VX_cyclic_arbiter.sv:32:9
			wire [NUM_REQS - 1:0] requests_w = (retain_grant ? prev_grant : requests);
			// Trace: src/VX_cyclic_arbiter.sv:33:9
			always @(posedge clk)
				// Trace: src/VX_cyclic_arbiter.sv:34:13
				if (reset)
					// Trace: src/VX_cyclic_arbiter.sv:35:17
					grant_index_r <= 1'sb0;
				else if ((grant_valid && grant_ready) && ~retain_grant) begin
					begin
						// Trace: src/VX_cyclic_arbiter.sv:37:17
						if (!IS_POW2 && (grant_index == sv2v_cast_76B5F_signed(NUM_REQS - 1)))
							// Trace: src/VX_cyclic_arbiter.sv:38:21
							grant_index_r <= 1'sb0;
						else
							// Trace: src/VX_cyclic_arbiter.sv:40:21
							grant_index_r <= grant_index + sv2v_cast_76B5F_signed(1);
					end
				end
			// Trace: src/VX_cyclic_arbiter.sv:44:9
			wire grant_valid_w;
			// Trace: src/VX_cyclic_arbiter.sv:45:9
			VX_priority_encoder #(.N(NUM_REQS)) grant_sel(
				.data_in(requests_w),
				.onehot_out(grant_onehot_um),
				.index_out(grant_index_um),
				.valid_out(grant_valid_w)
			);
			// Trace: src/VX_cyclic_arbiter.sv:53:9
			VX_demux #(
				.DATAW(1),
				.N(NUM_REQS)
			) grant_decoder(
				.sel_in(grant_index_r),
				.data_in(1'b1),
				.data_out(grant_onehot_w)
			);
			// Trace: src/VX_cyclic_arbiter.sv:61:9
			wire is_hit = requests[grant_index_r] && ~retain_grant;
			// Trace: src/VX_cyclic_arbiter.sv:62:9
			assign grant_index = (is_hit ? grant_index_r : grant_index_um);
			// Trace: src/VX_cyclic_arbiter.sv:63:9
			assign grant_onehot = (is_hit ? grant_onehot_w : grant_onehot_um);
			// Trace: src/VX_cyclic_arbiter.sv:64:9
			assign grant_valid = (STICKY != 0 ? |requests : grant_valid_w);
		end
	endgenerate
endmodule
// removed interface: VX_decode_if
// removed interface: VX_dcr_bus_if
module VX_fifo_queue (
	clk,
	reset,
	push,
	pop,
	data_in,
	data_out,
	empty,
	alm_empty,
	full,
	alm_full,
	size
);
	// Trace: src/VX_fifo_queue.sv:2:15
	parameter DATAW = 32;
	// Trace: src/VX_fifo_queue.sv:3:15
	parameter DEPTH = 32;
	// Trace: src/VX_fifo_queue.sv:4:15
	parameter ALM_FULL = DEPTH - 1;
	// Trace: src/VX_fifo_queue.sv:5:15
	parameter ALM_EMPTY = 1;
	// Trace: src/VX_fifo_queue.sv:6:15
	parameter OUT_REG = 0;
	// Trace: src/VX_fifo_queue.sv:7:15
	parameter LUTRAM = 0;
	// Trace: src/VX_fifo_queue.sv:8:15
	parameter SIZEW = $clog2(DEPTH + 1);
	// Trace: src/VX_fifo_queue.sv:10:5
	input wire clk;
	// Trace: src/VX_fifo_queue.sv:11:5
	input wire reset;
	// Trace: src/VX_fifo_queue.sv:12:5
	input wire push;
	// Trace: src/VX_fifo_queue.sv:13:5
	input wire pop;
	// Trace: src/VX_fifo_queue.sv:14:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_fifo_queue.sv:15:5
	output wire [DATAW - 1:0] data_out;
	// Trace: src/VX_fifo_queue.sv:16:5
	output wire empty;
	// Trace: src/VX_fifo_queue.sv:17:5
	output wire alm_empty;
	// Trace: src/VX_fifo_queue.sv:18:5
	output wire full;
	// Trace: src/VX_fifo_queue.sv:19:5
	output wire alm_full;
	// Trace: src/VX_fifo_queue.sv:20:5
	output wire [SIZEW - 1:0] size;
	// Trace: src/VX_fifo_queue.sv:22:5
	VX_pending_size #(
		.SIZE(DEPTH),
		.ALM_EMPTY(ALM_EMPTY),
		.ALM_FULL(ALM_FULL)
	) pending_size(
		.clk(clk),
		.reset(reset),
		.incr(push),
		.decr(pop),
		.empty(empty),
		.full(full),
		.alm_empty(alm_empty),
		.alm_full(alm_full),
		.size(size)
	);
	// Trace: src/VX_fifo_queue.sv:37:5
	generate
		if (DEPTH == 1) begin : g_depth_1
			// Trace: src/VX_fifo_queue.sv:38:9
			reg [DATAW - 1:0] head_r;
			// Trace: src/VX_fifo_queue.sv:39:9
			always @(posedge clk)
				// Trace: src/VX_fifo_queue.sv:40:13
				if (push)
					// Trace: src/VX_fifo_queue.sv:41:17
					head_r <= data_in;
			// Trace: src/VX_fifo_queue.sv:44:9
			assign data_out = head_r;
		end
		else begin : g_depth_n
			// Trace: src/VX_fifo_queue.sv:46:9
			localparam ADDRW = $clog2(DEPTH);
			// Trace: src/VX_fifo_queue.sv:47:9
			wire [DATAW - 1:0] data_out_w;
			// Trace: src/VX_fifo_queue.sv:48:9
			reg [ADDRW - 1:0] rd_ptr_r;
			// Trace: src/VX_fifo_queue.sv:49:9
			reg [ADDRW - 1:0] wr_ptr_r;
			// Trace: src/VX_fifo_queue.sv:50:9
			always @(posedge clk)
				// Trace: src/VX_fifo_queue.sv:51:13
				if (reset) begin
					// Trace: src/VX_fifo_queue.sv:52:17
					wr_ptr_r <= 1'sb0;
					// Trace: src/VX_fifo_queue.sv:53:17
					rd_ptr_r <= (OUT_REG != 0 ? 1 : 0);
				end
				else begin
					// Trace: src/VX_fifo_queue.sv:55:17
					begin : sv2v_autoblock_1
						reg [ADDRW - 1:0] sv2v_tmp_cast;
						sv2v_tmp_cast = push;
						wr_ptr_r <= wr_ptr_r + sv2v_tmp_cast;
					end
					// Trace: src/VX_fifo_queue.sv:56:17
					begin : sv2v_autoblock_2
						reg [ADDRW - 1:0] sv2v_tmp_cast_1;
						sv2v_tmp_cast_1 = pop;
						rd_ptr_r <= rd_ptr_r + sv2v_tmp_cast_1;
					end
				end
			// Trace: src/VX_fifo_queue.sv:59:9
			VX_dp_ram #(
				.DATAW(DATAW),
				.SIZE(DEPTH),
				.LUTRAM(LUTRAM),
				.RDW_MODE("W"),
				.RADDR_REG(1),
				.RADDR_RESET(1)
			) dp_ram(
				.clk(clk),
				.reset(reset),
				.read(1'b1),
				.write(push),
				.wren(1'b1),
				.raddr(rd_ptr_r),
				.waddr(wr_ptr_r),
				.wdata(data_in),
				.rdata(data_out_w)
			);
			if (OUT_REG != 0) begin : g_out_reg
				// Trace: src/VX_fifo_queue.sv:78:13
				reg [DATAW - 1:0] data_out_r;
				// Trace: src/VX_fifo_queue.sv:79:13
				function automatic signed [ADDRW - 1:0] sv2v_cast_8BB5D_signed;
					input reg signed [ADDRW - 1:0] inp;
					sv2v_cast_8BB5D_signed = inp;
				endfunction
				wire going_empty = (ALM_EMPTY == 1 ? alm_empty : size[ADDRW - 1:0] == sv2v_cast_8BB5D_signed(1));
				// Trace: src/VX_fifo_queue.sv:80:13
				wire bypass = push && (empty || (going_empty && pop));
				// Trace: src/VX_fifo_queue.sv:81:13
				always @(posedge clk)
					// Trace: src/VX_fifo_queue.sv:82:17
					if (bypass)
						// Trace: src/VX_fifo_queue.sv:83:21
						data_out_r <= data_in;
					else if (pop)
						// Trace: src/VX_fifo_queue.sv:85:21
						data_out_r <= data_out_w;
				// Trace: src/VX_fifo_queue.sv:88:13
				assign data_out = data_out_r;
			end
			else begin : g_no_out_reg
				// Trace: src/VX_fifo_queue.sv:90:13
				assign data_out = data_out_w;
			end
		end
	endgenerate
endmodule
module VX_generic_arbiter (
	clk,
	reset,
	requests,
	grant_index,
	grant_onehot,
	grant_valid,
	grant_ready
);
	// Trace: src/VX_generic_arbiter.sv:2:15
	parameter NUM_REQS = 1;
	// Trace: src/VX_generic_arbiter.sv:3:15
	parameter TYPE = "P";
	// Trace: src/VX_generic_arbiter.sv:4:15
	parameter STICKY = 0;
	// Trace: src/VX_generic_arbiter.sv:5:15
	parameter LOG_NUM_REQS = (NUM_REQS > 1 ? $clog2(NUM_REQS) : 1);
	// Trace: src/VX_generic_arbiter.sv:7:5
	input wire clk;
	// Trace: src/VX_generic_arbiter.sv:8:5
	input wire reset;
	// Trace: src/VX_generic_arbiter.sv:9:5
	input wire [NUM_REQS - 1:0] requests;
	// Trace: src/VX_generic_arbiter.sv:10:5
	output wire [LOG_NUM_REQS - 1:0] grant_index;
	// Trace: src/VX_generic_arbiter.sv:11:5
	output wire [NUM_REQS - 1:0] grant_onehot;
	// Trace: src/VX_generic_arbiter.sv:12:5
	output wire grant_valid;
	// Trace: src/VX_generic_arbiter.sv:13:5
	input wire grant_ready;
	// Trace: src/VX_generic_arbiter.sv:15:5
	generate
		if (TYPE == "P") begin : g_priority
			// Trace: src/VX_generic_arbiter.sv:16:9
			VX_priority_arbiter #(
				.NUM_REQS(NUM_REQS),
				.STICKY(STICKY)
			) priority_arbiter(
				.clk(clk),
				.reset(reset),
				.requests(requests),
				.grant_valid(grant_valid),
				.grant_index(grant_index),
				.grant_onehot(grant_onehot),
				.grant_ready(grant_ready)
			);
		end
		else if (TYPE == "R") begin : g_round_robin
			// Trace: src/VX_generic_arbiter.sv:29:9
			VX_rr_arbiter #(
				.NUM_REQS(NUM_REQS),
				.STICKY(STICKY)
			) rr_arbiter(
				.clk(clk),
				.reset(reset),
				.requests(requests),
				.grant_valid(grant_valid),
				.grant_index(grant_index),
				.grant_onehot(grant_onehot),
				.grant_ready(grant_ready)
			);
		end
		else if (TYPE == "M") begin : g_matrix
			// Trace: src/VX_generic_arbiter.sv:42:9
			VX_matrix_arbiter #(
				.NUM_REQS(NUM_REQS),
				.STICKY(STICKY)
			) matrix_arbiter(
				.clk(clk),
				.reset(reset),
				.requests(requests),
				.grant_valid(grant_valid),
				.grant_index(grant_index),
				.grant_onehot(grant_onehot),
				.grant_ready(grant_ready)
			);
		end
		else if (TYPE == "C") begin : g_cyclic
			// Trace: src/VX_generic_arbiter.sv:55:9
			VX_cyclic_arbiter #(
				.NUM_REQS(NUM_REQS),
				.STICKY(STICKY)
			) cyclic_arbiter(
				.clk(clk),
				.reset(reset),
				.requests(requests),
				.grant_valid(grant_valid),
				.grant_index(grant_index),
				.grant_onehot(grant_onehot),
				.grant_ready(grant_ready)
			);
		end
	endgenerate
endmodule
// removed package "VX_fpu_pkg"
// removed module with interface ports: VX_dcr_data
module VX_shift_register (
	clk,
	reset,
	enable,
	data_in,
	data_out
);
	// Trace: src/VX_shift_register.sv:2:15
	parameter DATAW = 1;
	// Trace: src/VX_shift_register.sv:3:15
	parameter RESETW = 0;
	// Trace: src/VX_shift_register.sv:4:15
	parameter DEPTH = 1;
	// Trace: src/VX_shift_register.sv:5:15
	parameter NUM_TAPS = 1;
	// Trace: src/VX_shift_register.sv:6:15
	parameter TAP_START = DEPTH - 1;
	// Trace: src/VX_shift_register.sv:7:15
	parameter TAP_STRIDE = 1;
	// Trace: src/VX_shift_register.sv:8:15
	parameter [(RESETW > 0 ? RESETW : 1) - 1:0] INIT_VALUE = {(RESETW > 0 ? RESETW : 1) {1'b0}};
	// Trace: src/VX_shift_register.sv:10:5
	input wire clk;
	// Trace: src/VX_shift_register.sv:11:5
	input wire reset;
	// Trace: src/VX_shift_register.sv:12:5
	input wire enable;
	// Trace: src/VX_shift_register.sv:13:5
	input wire [DATAW - 1:0] data_in;
	// Trace: src/VX_shift_register.sv:14:5
	output wire [(NUM_TAPS * DATAW) - 1:0] data_out;
	// Trace: src/VX_shift_register.sv:17:5
	generate
		if (DEPTH == 0) begin : g_passthru
			// Trace: src/VX_shift_register.sv:18:9
			assign data_out = data_in;
		end
		else begin : g_shift
			// Trace: src/VX_shift_register.sv:20:9
			reg [(DEPTH * DATAW) - 1:0] pipe;
			if (RESETW == DATAW) begin : g_full_reset
				genvar _gv_i_209;
				for (_gv_i_209 = 0; _gv_i_209 < DEPTH; _gv_i_209 = _gv_i_209 + 1) begin : g_stages
					localparam i = _gv_i_209;
					// Trace: src/VX_shift_register.sv:23:17
					always @(posedge clk)
						// Trace: src/VX_shift_register.sv:24:21
						if (reset)
							// Trace: src/VX_shift_register.sv:25:25
							pipe[i * DATAW+:DATAW] <= INIT_VALUE;
						else if (enable)
							// Trace: src/VX_shift_register.sv:27:25
							pipe[i * DATAW+:DATAW] <= (i == 0 ? data_in : pipe[(i - 1) * DATAW+:DATAW]);
				end
			end
			else if (RESETW != 0) begin : g_partial_reset
				genvar _gv_i_210;
				for (_gv_i_210 = 0; _gv_i_210 < DEPTH; _gv_i_210 = _gv_i_210 + 1) begin : g_stages
					localparam i = _gv_i_210;
					// Trace: src/VX_shift_register.sv:33:17
					always @(posedge clk)
						// Trace: src/VX_shift_register.sv:34:21
						if (reset)
							// Trace: src/VX_shift_register.sv:35:25
							pipe[(i * DATAW) + ((DATAW - 1) >= (DATAW - RESETW) ? DATAW - 1 : ((DATAW - 1) + ((DATAW - 1) >= (DATAW - RESETW) ? ((DATAW - 1) - (DATAW - RESETW)) + 1 : ((DATAW - RESETW) - (DATAW - 1)) + 1)) - 1)-:((DATAW - 1) >= (DATAW - RESETW) ? ((DATAW - 1) - (DATAW - RESETW)) + 1 : ((DATAW - RESETW) - (DATAW - 1)) + 1)] <= INIT_VALUE;
						else if (enable)
							// Trace: src/VX_shift_register.sv:37:25
							pipe[(i * DATAW) + ((DATAW - 1) >= (DATAW - RESETW) ? DATAW - 1 : ((DATAW - 1) + ((DATAW - 1) >= (DATAW - RESETW) ? ((DATAW - 1) - (DATAW - RESETW)) + 1 : ((DATAW - RESETW) - (DATAW - 1)) + 1)) - 1)-:((DATAW - 1) >= (DATAW - RESETW) ? ((DATAW - 1) - (DATAW - RESETW)) + 1 : ((DATAW - RESETW) - (DATAW - 1)) + 1)] <= (i == 0 ? data_in[DATAW - 1:DATAW - RESETW] : pipe[((i - 1) * DATAW) + ((DATAW - 1) >= (DATAW - RESETW) ? DATAW - 1 : ((DATAW - 1) + ((DATAW - 1) >= (DATAW - RESETW) ? ((DATAW - 1) - (DATAW - RESETW)) + 1 : ((DATAW - RESETW) - (DATAW - 1)) + 1)) - 1)-:((DATAW - 1) >= (DATAW - RESETW) ? ((DATAW - 1) - (DATAW - RESETW)) + 1 : ((DATAW - RESETW) - (DATAW - 1)) + 1)]);
					// Trace: src/VX_shift_register.sv:40:17
					always @(posedge clk)
						// Trace: src/VX_shift_register.sv:41:21
						if (enable)
							// Trace: src/VX_shift_register.sv:42:25
							pipe[(i * DATAW) + ((DATAW - RESETW) - 1)-:DATAW - RESETW] <= (i == 0 ? data_in[(DATAW - RESETW) - 1:0] : pipe[((i - 1) * DATAW) + ((DATAW - RESETW) - 1)-:DATAW - RESETW]);
				end
			end
			else begin : g_no_reset
				genvar _gv_i_211;
				for (_gv_i_211 = 0; _gv_i_211 < DEPTH; _gv_i_211 = _gv_i_211 + 1) begin : g_stages
					localparam i = _gv_i_211;
					// Trace: src/VX_shift_register.sv:48:17
					always @(posedge clk)
						// Trace: src/VX_shift_register.sv:49:21
						if (enable)
							// Trace: src/VX_shift_register.sv:50:25
							pipe[i * DATAW+:DATAW] <= (i == 0 ? data_in : pipe[(i - 1) * DATAW+:DATAW]);
				end
			end
			genvar _gv_i_212;
			for (_gv_i_212 = 0; _gv_i_212 < NUM_TAPS; _gv_i_212 = _gv_i_212 + 1) begin : g_taps
				localparam i = _gv_i_212;
				// Trace: src/VX_shift_register.sv:56:13
				assign data_out[i * DATAW+:DATAW] = pipe[((i * TAP_STRIDE) + TAP_START) * DATAW+:DATAW];
			end
		end
	endgenerate
endmodule
module VX_lzc (
	data_in,
	data_out,
	valid_out
);
	// Trace: src/VX_lzc.sv:2:15
	parameter N = 2;
	// Trace: src/VX_lzc.sv:3:15
	parameter REVERSE = 0;
	// Trace: src/VX_lzc.sv:4:15
	parameter LOGN = (N > 1 ? $clog2(N) : 1);
	// Trace: src/VX_lzc.sv:6:5
	input wire [N - 1:0] data_in;
	// Trace: src/VX_lzc.sv:7:5
	output wire [LOGN - 1:0] data_out;
	// Trace: src/VX_lzc.sv:8:5
	output wire valid_out;
	// Trace: src/VX_lzc.sv:10:5
	function automatic signed [LOGN - 1:0] sv2v_cast_B9644_signed;
		input reg signed [LOGN - 1:0] inp;
		sv2v_cast_B9644_signed = inp;
	endfunction
	generate
		if (N == 1) begin : g_passthru
			// Trace: src/VX_lzc.sv:11:9
			assign data_out = 1'sb0;
			// Trace: src/VX_lzc.sv:12:9
			assign valid_out = data_in;
		end
		else begin : g_lzc
			// Trace: src/VX_lzc.sv:14:9
			wire [(N * LOGN) - 1:0] indices;
			genvar _gv_i_213;
			for (_gv_i_213 = 0; _gv_i_213 < N; _gv_i_213 = _gv_i_213 + 1) begin : g_indices
				localparam i = _gv_i_213;
				// Trace: src/VX_lzc.sv:16:13
				assign indices[i * LOGN+:LOGN] = (REVERSE ? sv2v_cast_B9644_signed(i) : sv2v_cast_B9644_signed((N - 1) - i));
			end
			// Trace: src/VX_lzc.sv:18:9
			VX_find_first #(
				.N(N),
				.DATAW(LOGN),
				.REVERSE(!REVERSE)
			) find_first(
				.valid_in(data_in),
				.data_in(indices),
				.data_out(data_out),
				.valid_out(valid_out)
			);
		end
	endgenerate
endmodule
module VX_multiplier (
	clk,
	enable,
	dataa,
	datab,
	result
);
	// Trace: src/VX_multiplier.sv:2:15
	parameter A_WIDTH = 1;
	// Trace: src/VX_multiplier.sv:3:15
	parameter B_WIDTH = A_WIDTH;
	// Trace: src/VX_multiplier.sv:4:15
	parameter R_WIDTH = A_WIDTH + B_WIDTH;
	// Trace: src/VX_multiplier.sv:5:15
	parameter SIGNED = 0;
	// Trace: src/VX_multiplier.sv:6:15
	parameter LATENCY = 0;
	// Trace: src/VX_multiplier.sv:8:5
	input wire clk;
	// Trace: src/VX_multiplier.sv:9:5
	input wire enable;
	// Trace: src/VX_multiplier.sv:10:5
	input wire [A_WIDTH - 1:0] dataa;
	// Trace: src/VX_multiplier.sv:11:5
	input wire [B_WIDTH - 1:0] datab;
	// Trace: src/VX_multiplier.sv:12:5
	output wire [R_WIDTH - 1:0] result;
	// Trace: src/VX_multiplier.sv:14:5
	wire [R_WIDTH - 1:0] prod_w;
	// Trace: src/VX_multiplier.sv:15:5
	function automatic [R_WIDTH - 1:0] sv2v_cast_875D6;
		input reg [R_WIDTH - 1:0] inp;
		sv2v_cast_875D6 = inp;
	endfunction
	function automatic signed [R_WIDTH - 1:0] sv2v_cast_875D6_signed;
		input reg signed [R_WIDTH - 1:0] inp;
		sv2v_cast_875D6_signed = inp;
	endfunction
	generate
		if (SIGNED != 0) begin : g_prod_s
			// Trace: src/VX_multiplier.sv:16:9
			assign prod_w = sv2v_cast_875D6_signed($signed(dataa) * $signed(datab));
		end
		else begin : g_prod_u
			// Trace: src/VX_multiplier.sv:18:9
			assign prod_w = sv2v_cast_875D6(dataa * datab);
		end
	endgenerate
	// Trace: src/VX_multiplier.sv:20:5
	VX_pipe_register #(
		.DATAW(R_WIDTH),
		.DEPTH(LATENCY)
	) pipe_reg(
		.clk(clk),
		.enable(enable),
		.reset(1'b0),
		.data_in(prod_w),
		.data_out(result)
	);
endmodule
// removed interface: VX_lsu_mem_if
// removed package "VX_gpu_pkg"
// removed module with interface ports: VX_cache_init
// removed interface: VX_decode_sched_if
// removed interface: VX_branch_ctl_if
module VX_elastic_adapter (
	clk,
	reset,
	valid_in,
	ready_in,
	ready_out,
	valid_out,
	busy,
	strobe
);
	// Trace: src/VX_elastic_adapter.sv:2:5
	input wire clk;
	// Trace: src/VX_elastic_adapter.sv:3:5
	input wire reset;
	// Trace: src/VX_elastic_adapter.sv:4:5
	input wire valid_in;
	// Trace: src/VX_elastic_adapter.sv:5:5
	output wire ready_in;
	// Trace: src/VX_elastic_adapter.sv:6:5
	input wire ready_out;
	// Trace: src/VX_elastic_adapter.sv:7:5
	output wire valid_out;
	// Trace: src/VX_elastic_adapter.sv:8:5
	input wire busy;
	// Trace: src/VX_elastic_adapter.sv:9:5
	output wire strobe;
	// Trace: src/VX_elastic_adapter.sv:11:5
	wire push = valid_in && ready_in;
	// Trace: src/VX_elastic_adapter.sv:12:5
	wire pop = valid_out && ready_out;
	// Trace: src/VX_elastic_adapter.sv:13:5
	reg loaded;
	// Trace: src/VX_elastic_adapter.sv:14:5
	always @(posedge clk)
		// Trace: src/VX_elastic_adapter.sv:15:9
		if (reset)
			// Trace: src/VX_elastic_adapter.sv:16:13
			loaded <= 0;
		else begin
			// Trace: src/VX_elastic_adapter.sv:18:13
			if (push)
				// Trace: src/VX_elastic_adapter.sv:19:17
				loaded <= 1;
			if (pop)
				// Trace: src/VX_elastic_adapter.sv:22:17
				loaded <= 0;
		end
	// Trace: src/VX_elastic_adapter.sv:26:5
	assign ready_in = ~loaded;
	// Trace: src/VX_elastic_adapter.sv:27:5
	assign valid_out = loaded && ~busy;
	// Trace: src/VX_elastic_adapter.sv:28:5
	assign strobe = push;
endmodule
// removed module with interface ports: VX_csr_data
// removed module with interface ports: VX_gbar_unit
// removed module with interface ports: VX_cache
// removed module with interface ports: VX_uop_sequencer
module VX_reset_relay (
	clk,
	reset,
	reset_o
);
	// Trace: src/VX_reset_relay.sv:2:15
	parameter N = 1;
	// Trace: src/VX_reset_relay.sv:3:15
	parameter MAX_FANOUT = 0;
	// Trace: src/VX_reset_relay.sv:5:5
	input wire clk;
	// Trace: src/VX_reset_relay.sv:6:5
	input wire reset;
	// Trace: src/VX_reset_relay.sv:7:5
	output wire [N - 1:0] reset_o;
	// Trace: src/VX_reset_relay.sv:9:5
	generate
		if ((MAX_FANOUT >= 0) && (N > (MAX_FANOUT + (MAX_FANOUT / 2)))) begin : g_relay
			// Trace: src/VX_reset_relay.sv:10:9
			localparam F = (MAX_FANOUT > 0 ? MAX_FANOUT : 1);
			// Trace: src/VX_reset_relay.sv:11:9
			localparam R = N / F;
			// Trace: src/VX_reset_relay.sv:12:10
			reg [R - 1:0] reset_r;
			genvar _gv_i_244;
			for (_gv_i_244 = 0; _gv_i_244 < R; _gv_i_244 = _gv_i_244 + 1) begin : g_reset_r
				localparam i = _gv_i_244;
				// Trace: src/VX_reset_relay.sv:14:13
				always @(posedge clk)
					// Trace: src/VX_reset_relay.sv:15:17
					reset_r[i] <= reset;
			end
			genvar _gv_i_245;
			for (_gv_i_245 = 0; _gv_i_245 < N; _gv_i_245 = _gv_i_245 + 1) begin : g_reset_o
				localparam i = _gv_i_245;
				// Trace: src/VX_reset_relay.sv:19:13
				assign reset_o[i] = reset_r[i / F];
			end
		end
		else begin : g_passthru
			// Trace: src/VX_reset_relay.sv:22:9
			assign reset_o = {N {reset}};
		end
	endgenerate
endmodule
// removed interface: VX_fpu_csr_if
// removed module with interface ports: VX_cluster
// removed interface: VX_mem_bus_if